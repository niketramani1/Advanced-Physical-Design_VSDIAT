magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1260 -1320 9135 51880
<< locali >>
rect 4744 50462 4760 50496
rect 4794 50462 5963 50496
rect 7280 50423 7857 50457
rect 5064 50350 5080 50384
rect 5114 50350 5853 50384
rect 5704 50260 5720 50294
rect 5754 50260 5963 50294
rect 5704 50036 5720 50070
rect 5754 50036 5963 50070
rect 5064 49946 5080 49980
rect 5114 49946 5853 49980
rect 7280 49873 7857 49907
rect 4664 49834 4680 49868
rect 4714 49834 5963 49868
rect 4584 49672 4600 49706
rect 4634 49672 5963 49706
rect 7280 49633 7857 49667
rect 5064 49560 5080 49594
rect 5114 49560 5853 49594
rect 5704 49470 5720 49504
rect 5754 49470 5963 49504
rect 5704 49246 5720 49280
rect 5754 49246 5963 49280
rect 5064 49156 5080 49190
rect 5114 49156 5853 49190
rect 7280 49083 7857 49117
rect 4504 49044 4520 49078
rect 4554 49044 5963 49078
rect 4744 48882 4760 48916
rect 4794 48882 5963 48916
rect 7280 48843 7857 48877
rect 4984 48770 5000 48804
rect 5034 48770 5853 48804
rect 5704 48680 5720 48714
rect 5754 48680 5963 48714
rect 5704 48456 5720 48490
rect 5754 48456 5963 48490
rect 4984 48366 5000 48400
rect 5034 48366 5853 48400
rect 7280 48293 7857 48327
rect 4664 48254 4680 48288
rect 4714 48254 5963 48288
rect 4584 48092 4600 48126
rect 4634 48092 5963 48126
rect 7280 48053 7857 48087
rect 4984 47980 5000 48014
rect 5034 47980 5853 48014
rect 5704 47890 5720 47924
rect 5754 47890 5963 47924
rect 5704 47666 5720 47700
rect 5754 47666 5963 47700
rect 4984 47576 5000 47610
rect 5034 47576 5853 47610
rect 7280 47503 7857 47537
rect 4504 47464 4520 47498
rect 4554 47464 5963 47498
rect 4744 47302 4760 47336
rect 4794 47302 5963 47336
rect 7280 47263 7857 47297
rect 4904 47190 4920 47224
rect 4954 47190 5853 47224
rect 5704 47100 5720 47134
rect 5754 47100 5963 47134
rect 5704 46876 5720 46910
rect 5754 46876 5963 46910
rect 4904 46786 4920 46820
rect 4954 46786 5853 46820
rect 7280 46713 7857 46747
rect 4664 46674 4680 46708
rect 4714 46674 5963 46708
rect 4584 46512 4600 46546
rect 4634 46512 5963 46546
rect 7280 46473 7857 46507
rect 4904 46400 4920 46434
rect 4954 46400 5853 46434
rect 5704 46310 5720 46344
rect 5754 46310 5963 46344
rect 5704 46086 5720 46120
rect 5754 46086 5963 46120
rect 4904 45996 4920 46030
rect 4954 45996 5853 46030
rect 7280 45923 7857 45957
rect 4504 45884 4520 45918
rect 4554 45884 5963 45918
rect 4744 45722 4760 45756
rect 4794 45722 5963 45756
rect 7280 45683 7857 45717
rect 4824 45610 4840 45644
rect 4874 45610 5853 45644
rect 5704 45520 5720 45554
rect 5754 45520 5963 45554
rect 5704 45296 5720 45330
rect 5754 45296 5963 45330
rect 4824 45206 4840 45240
rect 4874 45206 5853 45240
rect 7280 45133 7857 45167
rect 4664 45094 4680 45128
rect 4714 45094 5963 45128
rect 4584 44932 4600 44966
rect 4634 44932 5963 44966
rect 7280 44893 7857 44927
rect 4824 44820 4840 44854
rect 4874 44820 5853 44854
rect 5704 44730 5720 44764
rect 5754 44730 5963 44764
rect 5704 44506 5720 44540
rect 5754 44506 5963 44540
rect 4824 44416 4840 44450
rect 4874 44416 5853 44450
rect 7280 44343 7857 44377
rect 4504 44304 4520 44338
rect 4554 44304 5963 44338
rect 4744 44142 4760 44176
rect 4794 44142 5963 44176
rect 7280 44103 7857 44137
rect 5064 44030 5080 44064
rect 5114 44030 5853 44064
rect 5624 43940 5640 43974
rect 5674 43940 5963 43974
rect 5624 43716 5640 43750
rect 5674 43716 5963 43750
rect 5064 43626 5080 43660
rect 5114 43626 5853 43660
rect 7280 43553 7857 43587
rect 4664 43514 4680 43548
rect 4714 43514 5963 43548
rect 4584 43352 4600 43386
rect 4634 43352 5963 43386
rect 7280 43313 7857 43347
rect 5064 43240 5080 43274
rect 5114 43240 5853 43274
rect 5624 43150 5640 43184
rect 5674 43150 5963 43184
rect 5624 42926 5640 42960
rect 5674 42926 5963 42960
rect 5064 42836 5080 42870
rect 5114 42836 5853 42870
rect 7280 42763 7857 42797
rect 4504 42724 4520 42758
rect 4554 42724 5963 42758
rect 4744 42562 4760 42596
rect 4794 42562 5963 42596
rect 7280 42523 7857 42557
rect 4984 42450 5000 42484
rect 5034 42450 5853 42484
rect 5624 42360 5640 42394
rect 5674 42360 5963 42394
rect 5624 42136 5640 42170
rect 5674 42136 5963 42170
rect 4984 42046 5000 42080
rect 5034 42046 5853 42080
rect 7280 41973 7857 42007
rect 4664 41934 4680 41968
rect 4714 41934 5963 41968
rect 4584 41772 4600 41806
rect 4634 41772 5963 41806
rect 7280 41733 7857 41767
rect 4984 41660 5000 41694
rect 5034 41660 5853 41694
rect 5624 41570 5640 41604
rect 5674 41570 5963 41604
rect 5624 41346 5640 41380
rect 5674 41346 5963 41380
rect 4984 41256 5000 41290
rect 5034 41256 5853 41290
rect 7280 41183 7857 41217
rect 4504 41144 4520 41178
rect 4554 41144 5963 41178
rect 4744 40982 4760 41016
rect 4794 40982 5963 41016
rect 7280 40943 7857 40977
rect 4904 40870 4920 40904
rect 4954 40870 5853 40904
rect 5624 40780 5640 40814
rect 5674 40780 5963 40814
rect 5624 40556 5640 40590
rect 5674 40556 5963 40590
rect 4904 40466 4920 40500
rect 4954 40466 5853 40500
rect 7280 40393 7857 40427
rect 4664 40354 4680 40388
rect 4714 40354 5963 40388
rect 4584 40192 4600 40226
rect 4634 40192 5963 40226
rect 7280 40153 7857 40187
rect 4904 40080 4920 40114
rect 4954 40080 5853 40114
rect 5624 39990 5640 40024
rect 5674 39990 5963 40024
rect 5624 39766 5640 39800
rect 5674 39766 5963 39800
rect 4904 39676 4920 39710
rect 4954 39676 5853 39710
rect 7280 39603 7857 39637
rect 4504 39564 4520 39598
rect 4554 39564 5963 39598
rect 4744 39402 4760 39436
rect 4794 39402 5963 39436
rect 7280 39363 7857 39397
rect 4824 39290 4840 39324
rect 4874 39290 5853 39324
rect 5624 39200 5640 39234
rect 5674 39200 5963 39234
rect 5624 38976 5640 39010
rect 5674 38976 5963 39010
rect 4824 38886 4840 38920
rect 4874 38886 5853 38920
rect 7280 38813 7857 38847
rect 4664 38774 4680 38808
rect 4714 38774 5963 38808
rect 4584 38612 4600 38646
rect 4634 38612 5963 38646
rect 7280 38573 7857 38607
rect 4824 38500 4840 38534
rect 4874 38500 5853 38534
rect 5624 38410 5640 38444
rect 5674 38410 5963 38444
rect 5624 38186 5640 38220
rect 5674 38186 5963 38220
rect 4824 38096 4840 38130
rect 4874 38096 5853 38130
rect 7280 38023 7857 38057
rect 4504 37984 4520 38018
rect 4554 37984 5963 38018
rect 4744 37822 4760 37856
rect 4794 37822 5963 37856
rect 7280 37783 7857 37817
rect 5064 37710 5080 37744
rect 5114 37710 5853 37744
rect 5544 37620 5560 37654
rect 5594 37620 5963 37654
rect 5544 37396 5560 37430
rect 5594 37396 5963 37430
rect 5064 37306 5080 37340
rect 5114 37306 5853 37340
rect 7280 37233 7857 37267
rect 4664 37194 4680 37228
rect 4714 37194 5963 37228
rect 4584 37032 4600 37066
rect 4634 37032 5963 37066
rect 7280 36993 7857 37027
rect 5064 36920 5080 36954
rect 5114 36920 5853 36954
rect 5544 36830 5560 36864
rect 5594 36830 5963 36864
rect 5544 36606 5560 36640
rect 5594 36606 5963 36640
rect 5064 36516 5080 36550
rect 5114 36516 5853 36550
rect 7280 36443 7857 36477
rect 4504 36404 4520 36438
rect 4554 36404 5963 36438
rect 4744 36242 4760 36276
rect 4794 36242 5963 36276
rect 7280 36203 7857 36237
rect 4984 36130 5000 36164
rect 5034 36130 5853 36164
rect 5544 36040 5560 36074
rect 5594 36040 5963 36074
rect 5544 35816 5560 35850
rect 5594 35816 5963 35850
rect 4984 35726 5000 35760
rect 5034 35726 5853 35760
rect 7280 35653 7857 35687
rect 4664 35614 4680 35648
rect 4714 35614 5963 35648
rect 4584 35452 4600 35486
rect 4634 35452 5963 35486
rect 7280 35413 7857 35447
rect 4984 35340 5000 35374
rect 5034 35340 5853 35374
rect 5544 35250 5560 35284
rect 5594 35250 5963 35284
rect 5544 35026 5560 35060
rect 5594 35026 5963 35060
rect 4984 34936 5000 34970
rect 5034 34936 5853 34970
rect 7280 34863 7857 34897
rect 4504 34824 4520 34858
rect 4554 34824 5963 34858
rect 4744 34662 4760 34696
rect 4794 34662 5963 34696
rect 7280 34623 7857 34657
rect 4904 34550 4920 34584
rect 4954 34550 5853 34584
rect 5544 34460 5560 34494
rect 5594 34460 5963 34494
rect 5544 34236 5560 34270
rect 5594 34236 5963 34270
rect 4904 34146 4920 34180
rect 4954 34146 5853 34180
rect 7280 34073 7857 34107
rect 4664 34034 4680 34068
rect 4714 34034 5963 34068
rect 4584 33872 4600 33906
rect 4634 33872 5963 33906
rect 7280 33833 7857 33867
rect 4904 33760 4920 33794
rect 4954 33760 5853 33794
rect 5544 33670 5560 33704
rect 5594 33670 5963 33704
rect 5544 33446 5560 33480
rect 5594 33446 5963 33480
rect 4904 33356 4920 33390
rect 4954 33356 5853 33390
rect 7280 33283 7857 33317
rect 4504 33244 4520 33278
rect 4554 33244 5963 33278
rect 4744 33082 4760 33116
rect 4794 33082 5963 33116
rect 7280 33043 7857 33077
rect 4824 32970 4840 33004
rect 4874 32970 5853 33004
rect 5544 32880 5560 32914
rect 5594 32880 5963 32914
rect 5544 32656 5560 32690
rect 5594 32656 5963 32690
rect 4824 32566 4840 32600
rect 4874 32566 5853 32600
rect 7280 32493 7857 32527
rect 4664 32454 4680 32488
rect 4714 32454 5963 32488
rect 4584 32292 4600 32326
rect 4634 32292 5963 32326
rect 7280 32253 7857 32287
rect 4824 32180 4840 32214
rect 4874 32180 5853 32214
rect 5544 32090 5560 32124
rect 5594 32090 5963 32124
rect 5544 31866 5560 31900
rect 5594 31866 5963 31900
rect 4824 31776 4840 31810
rect 4874 31776 5853 31810
rect 7280 31703 7857 31737
rect 4504 31664 4520 31698
rect 4554 31664 5963 31698
rect 4744 31502 4760 31536
rect 4794 31502 5963 31536
rect 7280 31463 7857 31497
rect 5064 31390 5080 31424
rect 5114 31390 5853 31424
rect 5464 31300 5480 31334
rect 5514 31300 5963 31334
rect 5464 31076 5480 31110
rect 5514 31076 5963 31110
rect 5064 30986 5080 31020
rect 5114 30986 5853 31020
rect 7280 30913 7857 30947
rect 4664 30874 4680 30908
rect 4714 30874 5963 30908
rect 4584 30712 4600 30746
rect 4634 30712 5963 30746
rect 7280 30673 7857 30707
rect 5064 30600 5080 30634
rect 5114 30600 5853 30634
rect 5464 30510 5480 30544
rect 5514 30510 5963 30544
rect 5464 30286 5480 30320
rect 5514 30286 5963 30320
rect 5064 30196 5080 30230
rect 5114 30196 5853 30230
rect 7280 30123 7857 30157
rect 4504 30084 4520 30118
rect 4554 30084 5963 30118
rect 4744 29922 4760 29956
rect 4794 29922 5963 29956
rect 7280 29883 7857 29917
rect 4984 29810 5000 29844
rect 5034 29810 5853 29844
rect 5464 29720 5480 29754
rect 5514 29720 5963 29754
rect 5464 29496 5480 29530
rect 5514 29496 5963 29530
rect 4984 29406 5000 29440
rect 5034 29406 5853 29440
rect 7280 29333 7857 29367
rect 4664 29294 4680 29328
rect 4714 29294 5963 29328
rect 4584 29132 4600 29166
rect 4634 29132 5963 29166
rect 7280 29093 7857 29127
rect 4984 29020 5000 29054
rect 5034 29020 5853 29054
rect 5464 28930 5480 28964
rect 5514 28930 5963 28964
rect 5464 28706 5480 28740
rect 5514 28706 5963 28740
rect 4984 28616 5000 28650
rect 5034 28616 5853 28650
rect 7280 28543 7857 28577
rect 4504 28504 4520 28538
rect 4554 28504 5963 28538
rect 4744 28342 4760 28376
rect 4794 28342 5963 28376
rect 7280 28303 7857 28337
rect 4904 28230 4920 28264
rect 4954 28230 5853 28264
rect 5464 28140 5480 28174
rect 5514 28140 5963 28174
rect 5464 27916 5480 27950
rect 5514 27916 5963 27950
rect 4904 27826 4920 27860
rect 4954 27826 5853 27860
rect 7280 27753 7857 27787
rect 4664 27714 4680 27748
rect 4714 27714 5963 27748
rect 4584 27552 4600 27586
rect 4634 27552 5963 27586
rect 7280 27513 7857 27547
rect 4904 27440 4920 27474
rect 4954 27440 5853 27474
rect 5464 27350 5480 27384
rect 5514 27350 5963 27384
rect 5464 27126 5480 27160
rect 5514 27126 5963 27160
rect 4904 27036 4920 27070
rect 4954 27036 5853 27070
rect 7280 26963 7857 26997
rect 4504 26924 4520 26958
rect 4554 26924 5963 26958
rect 4744 26762 4760 26796
rect 4794 26762 5963 26796
rect 7280 26723 7857 26757
rect 4824 26650 4840 26684
rect 4874 26650 5853 26684
rect 5464 26560 5480 26594
rect 5514 26560 5963 26594
rect 5464 26336 5480 26370
rect 5514 26336 5963 26370
rect 4824 26246 4840 26280
rect 4874 26246 5853 26280
rect 7280 26173 7857 26207
rect 4664 26134 4680 26168
rect 4714 26134 5963 26168
rect 4584 25972 4600 26006
rect 4634 25972 5963 26006
rect 7280 25933 7857 25967
rect 4824 25860 4840 25894
rect 4874 25860 5853 25894
rect 5464 25770 5480 25804
rect 5514 25770 5963 25804
rect 5464 25546 5480 25580
rect 5514 25546 5963 25580
rect 4824 25456 4840 25490
rect 4874 25456 5853 25490
rect 7280 25383 7857 25417
rect 4504 25344 4520 25378
rect 4554 25344 5963 25378
rect 4744 25182 4760 25216
rect 4794 25182 5963 25216
rect 7280 25143 7857 25177
rect 5064 25070 5080 25104
rect 5114 25070 5853 25104
rect 5384 24980 5400 25014
rect 5434 24980 5963 25014
rect 5384 24756 5400 24790
rect 5434 24756 5963 24790
rect 5064 24666 5080 24700
rect 5114 24666 5853 24700
rect 7280 24593 7857 24627
rect 4664 24554 4680 24588
rect 4714 24554 5963 24588
rect 4584 24392 4600 24426
rect 4634 24392 5963 24426
rect 7280 24353 7857 24387
rect 5064 24280 5080 24314
rect 5114 24280 5853 24314
rect 5384 24190 5400 24224
rect 5434 24190 5963 24224
rect 5384 23966 5400 24000
rect 5434 23966 5963 24000
rect 5064 23876 5080 23910
rect 5114 23876 5853 23910
rect 7280 23803 7857 23837
rect 4504 23764 4520 23798
rect 4554 23764 5963 23798
rect 4744 23602 4760 23636
rect 4794 23602 5963 23636
rect 7280 23563 7857 23597
rect 4984 23490 5000 23524
rect 5034 23490 5853 23524
rect 5384 23400 5400 23434
rect 5434 23400 5963 23434
rect 5384 23176 5400 23210
rect 5434 23176 5963 23210
rect 4984 23086 5000 23120
rect 5034 23086 5853 23120
rect 7280 23013 7857 23047
rect 4664 22974 4680 23008
rect 4714 22974 5963 23008
rect 4584 22812 4600 22846
rect 4634 22812 5963 22846
rect 7280 22773 7857 22807
rect 4984 22700 5000 22734
rect 5034 22700 5853 22734
rect 5384 22610 5400 22644
rect 5434 22610 5963 22644
rect 5384 22386 5400 22420
rect 5434 22386 5963 22420
rect 4984 22296 5000 22330
rect 5034 22296 5853 22330
rect 7280 22223 7857 22257
rect 4504 22184 4520 22218
rect 4554 22184 5963 22218
rect 4744 22022 4760 22056
rect 4794 22022 5963 22056
rect 7280 21983 7857 22017
rect 4904 21910 4920 21944
rect 4954 21910 5853 21944
rect 5384 21820 5400 21854
rect 5434 21820 5963 21854
rect 5384 21596 5400 21630
rect 5434 21596 5963 21630
rect 4904 21506 4920 21540
rect 4954 21506 5853 21540
rect 7280 21433 7857 21467
rect 4664 21394 4680 21428
rect 4714 21394 5963 21428
rect 4584 21232 4600 21266
rect 4634 21232 5963 21266
rect 7280 21193 7857 21227
rect 4904 21120 4920 21154
rect 4954 21120 5853 21154
rect 5384 21030 5400 21064
rect 5434 21030 5963 21064
rect 5384 20806 5400 20840
rect 5434 20806 5963 20840
rect 4904 20716 4920 20750
rect 4954 20716 5853 20750
rect 7280 20643 7857 20677
rect 4504 20604 4520 20638
rect 4554 20604 5963 20638
rect 4744 20442 4760 20476
rect 4794 20442 5963 20476
rect 7280 20403 7857 20437
rect 4824 20330 4840 20364
rect 4874 20330 5853 20364
rect 5384 20240 5400 20274
rect 5434 20240 5963 20274
rect 5384 20016 5400 20050
rect 5434 20016 5963 20050
rect 4824 19926 4840 19960
rect 4874 19926 5853 19960
rect 7280 19853 7857 19887
rect 4664 19814 4680 19848
rect 4714 19814 5963 19848
rect 4584 19652 4600 19686
rect 4634 19652 5963 19686
rect 7280 19613 7857 19647
rect 4824 19540 4840 19574
rect 4874 19540 5853 19574
rect 5384 19450 5400 19484
rect 5434 19450 5963 19484
rect 5384 19226 5400 19260
rect 5434 19226 5963 19260
rect 4824 19136 4840 19170
rect 4874 19136 5853 19170
rect 7280 19063 7857 19097
rect 4504 19024 4520 19058
rect 4554 19024 5963 19058
rect 4744 18862 4760 18896
rect 4794 18862 5963 18896
rect 7280 18823 7857 18857
rect 5064 18750 5080 18784
rect 5114 18750 5853 18784
rect 5304 18660 5320 18694
rect 5354 18660 5963 18694
rect 5304 18436 5320 18470
rect 5354 18436 5963 18470
rect 5064 18346 5080 18380
rect 5114 18346 5853 18380
rect 7280 18273 7857 18307
rect 4664 18234 4680 18268
rect 4714 18234 5963 18268
rect 4584 18072 4600 18106
rect 4634 18072 5963 18106
rect 7280 18033 7857 18067
rect 5064 17960 5080 17994
rect 5114 17960 5853 17994
rect 5304 17870 5320 17904
rect 5354 17870 5963 17904
rect 5304 17646 5320 17680
rect 5354 17646 5963 17680
rect 5064 17556 5080 17590
rect 5114 17556 5853 17590
rect 7280 17483 7857 17517
rect 4504 17444 4520 17478
rect 4554 17444 5963 17478
rect 4744 17282 4760 17316
rect 4794 17282 5963 17316
rect 7280 17243 7857 17277
rect 4984 17170 5000 17204
rect 5034 17170 5853 17204
rect 5304 17080 5320 17114
rect 5354 17080 5963 17114
rect 5304 16856 5320 16890
rect 5354 16856 5963 16890
rect 4984 16766 5000 16800
rect 5034 16766 5853 16800
rect 7280 16693 7857 16727
rect 4664 16654 4680 16688
rect 4714 16654 5963 16688
rect 4584 16492 4600 16526
rect 4634 16492 5963 16526
rect 7280 16453 7857 16487
rect 4984 16380 5000 16414
rect 5034 16380 5853 16414
rect 5304 16290 5320 16324
rect 5354 16290 5963 16324
rect 5304 16066 5320 16100
rect 5354 16066 5963 16100
rect 4984 15976 5000 16010
rect 5034 15976 5853 16010
rect 7280 15903 7857 15937
rect 4504 15864 4520 15898
rect 4554 15864 5963 15898
rect 4744 15702 4760 15736
rect 4794 15702 5963 15736
rect 7280 15663 7857 15697
rect 4904 15590 4920 15624
rect 4954 15590 5853 15624
rect 5304 15500 5320 15534
rect 5354 15500 5963 15534
rect 5304 15276 5320 15310
rect 5354 15276 5963 15310
rect 4904 15186 4920 15220
rect 4954 15186 5853 15220
rect 7280 15113 7857 15147
rect 4664 15074 4680 15108
rect 4714 15074 5963 15108
rect 4584 14912 4600 14946
rect 4634 14912 5963 14946
rect 7280 14873 7857 14907
rect 4904 14800 4920 14834
rect 4954 14800 5853 14834
rect 5304 14710 5320 14744
rect 5354 14710 5963 14744
rect 5304 14486 5320 14520
rect 5354 14486 5963 14520
rect 4904 14396 4920 14430
rect 4954 14396 5853 14430
rect 7280 14323 7857 14357
rect 4504 14284 4520 14318
rect 4554 14284 5963 14318
rect 4744 14122 4760 14156
rect 4794 14122 5963 14156
rect 7280 14083 7857 14117
rect 4824 14010 4840 14044
rect 4874 14010 5853 14044
rect 5304 13920 5320 13954
rect 5354 13920 5963 13954
rect 5304 13696 5320 13730
rect 5354 13696 5963 13730
rect 4824 13606 4840 13640
rect 4874 13606 5853 13640
rect 7280 13533 7857 13567
rect 4664 13494 4680 13528
rect 4714 13494 5963 13528
rect 4584 13332 4600 13366
rect 4634 13332 5963 13366
rect 7280 13293 7857 13327
rect 4824 13220 4840 13254
rect 4874 13220 5853 13254
rect 5304 13130 5320 13164
rect 5354 13130 5963 13164
rect 5304 12906 5320 12940
rect 5354 12906 5963 12940
rect 4824 12816 4840 12850
rect 4874 12816 5853 12850
rect 7280 12743 7857 12777
rect 4504 12704 4520 12738
rect 4554 12704 5963 12738
rect 4744 12542 4760 12576
rect 4794 12542 5963 12576
rect 7280 12503 7857 12537
rect 5064 12430 5080 12464
rect 5114 12430 5853 12464
rect 5224 12340 5240 12374
rect 5274 12340 5963 12374
rect 5224 12116 5240 12150
rect 5274 12116 5963 12150
rect 5064 12026 5080 12060
rect 5114 12026 5853 12060
rect 7280 11953 7857 11987
rect 4664 11914 4680 11948
rect 4714 11914 5963 11948
rect 4584 11752 4600 11786
rect 4634 11752 5963 11786
rect 7280 11713 7857 11747
rect 5064 11640 5080 11674
rect 5114 11640 5853 11674
rect 5224 11550 5240 11584
rect 5274 11550 5963 11584
rect 5224 11326 5240 11360
rect 5274 11326 5963 11360
rect 5064 11236 5080 11270
rect 5114 11236 5853 11270
rect 7280 11163 7857 11197
rect 4504 11124 4520 11158
rect 4554 11124 5963 11158
rect 4744 10962 4760 10996
rect 4794 10962 5963 10996
rect 7280 10923 7857 10957
rect 4984 10850 5000 10884
rect 5034 10850 5853 10884
rect 5224 10760 5240 10794
rect 5274 10760 5963 10794
rect 5224 10536 5240 10570
rect 5274 10536 5963 10570
rect 4984 10446 5000 10480
rect 5034 10446 5853 10480
rect 7280 10373 7857 10407
rect 4664 10334 4680 10368
rect 4714 10334 5963 10368
rect 4584 10172 4600 10206
rect 4634 10172 5963 10206
rect 7280 10133 7857 10167
rect 4984 10060 5000 10094
rect 5034 10060 5853 10094
rect 5224 9970 5240 10004
rect 5274 9970 5963 10004
rect 5224 9746 5240 9780
rect 5274 9746 5963 9780
rect 4984 9656 5000 9690
rect 5034 9656 5853 9690
rect 7280 9583 7857 9617
rect 4504 9544 4520 9578
rect 4554 9544 5963 9578
rect 4744 9382 4760 9416
rect 4794 9382 5963 9416
rect 7280 9343 7857 9377
rect 4904 9270 4920 9304
rect 4954 9270 5853 9304
rect 5224 9180 5240 9214
rect 5274 9180 5963 9214
rect 5224 8956 5240 8990
rect 5274 8956 5963 8990
rect 4904 8866 4920 8900
rect 4954 8866 5853 8900
rect 7280 8793 7857 8827
rect 4664 8754 4680 8788
rect 4714 8754 5963 8788
rect 4584 8592 4600 8626
rect 4634 8592 5963 8626
rect 7280 8553 7857 8587
rect 4904 8480 4920 8514
rect 4954 8480 5853 8514
rect 5224 8390 5240 8424
rect 5274 8390 5963 8424
rect 5224 8166 5240 8200
rect 5274 8166 5963 8200
rect 4904 8076 4920 8110
rect 4954 8076 5853 8110
rect 7280 8003 7857 8037
rect 4504 7964 4520 7998
rect 4554 7964 5963 7998
rect 4426 7797 4460 7813
rect 4744 7802 4760 7836
rect 4794 7802 5963 7836
rect 7280 7763 7857 7797
rect 4426 7747 4460 7763
rect 4824 7690 4840 7724
rect 4874 7690 5853 7724
rect 5224 7600 5240 7634
rect 5274 7600 5963 7634
rect 5224 7376 5240 7410
rect 5274 7376 5963 7410
rect 4824 7286 4840 7320
rect 4874 7286 5853 7320
rect 4426 7247 4460 7263
rect 7280 7213 7857 7247
rect 4426 7197 4460 7213
rect 4664 7174 4680 7208
rect 4714 7174 5963 7208
rect 4426 7007 4460 7023
rect 4584 7012 4600 7046
rect 4634 7012 5963 7046
rect 7280 6973 7857 7007
rect 4426 6957 4460 6973
rect 4824 6900 4840 6934
rect 4874 6900 5853 6934
rect 5224 6810 5240 6844
rect 5274 6810 5963 6844
rect 5224 6586 5240 6620
rect 5274 6586 5963 6620
rect 4824 6496 4840 6530
rect 4874 6496 5853 6530
rect 4426 6457 4460 6473
rect 7280 6423 7857 6457
rect 4426 6407 4460 6423
rect 4504 6384 4520 6418
rect 4554 6384 5963 6418
rect 4426 6217 4460 6233
rect 4744 6222 4760 6256
rect 4794 6222 5963 6256
rect 7280 6183 7857 6217
rect 4426 6167 4460 6183
rect 5064 6110 5080 6144
rect 5114 6110 5853 6144
rect 5144 6020 5160 6054
rect 5194 6020 5963 6054
rect 5144 5796 5160 5830
rect 5194 5796 5963 5830
rect 844 5717 878 5733
rect 480 5683 496 5717
rect 530 5683 844 5717
rect 5064 5706 5080 5740
rect 5114 5706 5853 5740
rect 844 5667 878 5683
rect 4426 5667 4460 5683
rect 7280 5633 7857 5667
rect 4426 5617 4460 5633
rect 4664 5594 4680 5628
rect 4714 5594 5963 5628
rect 4426 5427 4460 5443
rect 4584 5432 4600 5466
rect 4634 5432 5963 5466
rect 7280 5393 7857 5427
rect 764 5377 798 5393
rect 4426 5377 4460 5393
rect 400 5343 416 5377
rect 450 5343 764 5377
rect 764 5327 798 5343
rect 5064 5320 5080 5354
rect 5114 5320 5853 5354
rect 5144 5230 5160 5264
rect 5194 5230 5963 5264
rect 5144 5006 5160 5040
rect 5194 5006 5963 5040
rect 684 4927 718 4943
rect 320 4893 336 4927
rect 370 4893 684 4927
rect 5064 4916 5080 4950
rect 5114 4916 5853 4950
rect 684 4877 718 4893
rect 4426 4877 4460 4893
rect 7280 4843 7857 4877
rect 4426 4827 4460 4843
rect 4504 4804 4520 4838
rect 4554 4804 5963 4838
rect 4744 4642 4760 4676
rect 4794 4642 5963 4676
rect 7280 4603 7857 4637
rect 4984 4530 5000 4564
rect 5034 4530 5853 4564
rect 5144 4440 5160 4474
rect 5194 4440 5963 4474
rect 5144 4216 5160 4250
rect 5194 4216 5963 4250
rect 4984 4126 5000 4160
rect 5034 4126 5853 4160
rect 7280 4053 7857 4087
rect 4664 4014 4680 4048
rect 4714 4014 5963 4048
rect 4426 3847 4460 3863
rect 4584 3852 4600 3886
rect 4634 3852 5963 3886
rect 7280 3813 7857 3847
rect 4426 3797 4460 3813
rect 4984 3740 5000 3774
rect 5034 3740 5853 3774
rect 5144 3650 5160 3684
rect 5194 3650 5963 3684
rect 5144 3426 5160 3460
rect 5194 3426 5963 3460
rect 4984 3336 5000 3370
rect 5034 3336 5853 3370
rect 4426 3297 4460 3313
rect 7280 3263 7857 3297
rect 4426 3247 4460 3263
rect 4504 3224 4520 3258
rect 4554 3224 5963 3258
rect 4426 3057 4460 3073
rect 4744 3062 4760 3096
rect 4794 3062 5963 3096
rect 7280 3023 7857 3057
rect 1440 3007 1474 3023
rect 4426 3007 4460 3023
rect 240 2973 256 3007
rect 290 2973 1440 3007
rect 1440 2957 1474 2973
rect 4904 2950 4920 2984
rect 4954 2950 5853 2984
rect 5144 2860 5160 2894
rect 5194 2860 5963 2894
rect 5144 2636 5160 2670
rect 5194 2636 5963 2670
rect 1360 2557 1394 2573
rect 160 2523 176 2557
rect 210 2523 1360 2557
rect 4904 2546 4920 2580
rect 4954 2546 5853 2580
rect 1360 2507 1394 2523
rect 4426 2507 4460 2523
rect 7280 2473 7857 2507
rect 4426 2457 4460 2473
rect 4664 2434 4680 2468
rect 4714 2434 5963 2468
rect 4584 2272 4600 2306
rect 4634 2272 5963 2306
rect 7280 2233 7857 2267
rect 4904 2160 4920 2194
rect 4954 2160 5853 2194
rect 5144 2070 5160 2104
rect 5194 2070 5963 2104
rect 5144 1846 5160 1880
rect 5194 1846 5963 1880
rect 4904 1756 4920 1790
rect 4954 1756 5853 1790
rect 7280 1683 7857 1717
rect 4504 1644 4520 1678
rect 4554 1644 5963 1678
rect 4426 1477 4460 1493
rect 4744 1482 4760 1516
rect 4794 1482 5963 1516
rect 7280 1443 7857 1477
rect 4426 1427 4460 1443
rect 4824 1370 4840 1404
rect 4874 1370 5853 1404
rect 5144 1280 5160 1314
rect 5194 1280 5963 1314
rect 5144 1056 5160 1090
rect 5194 1056 5963 1090
rect 4824 966 4840 1000
rect 4874 966 5853 1000
rect 4426 927 4460 943
rect 7280 893 7857 927
rect 4426 877 4460 893
rect 4664 854 4680 888
rect 4714 854 5963 888
rect 4426 687 4460 703
rect 4584 692 4600 726
rect 4634 692 5963 726
rect 7280 653 7857 687
rect 1440 637 1474 653
rect 4426 637 4460 653
rect 80 603 96 637
rect 130 603 1440 637
rect 1440 587 1474 603
rect 4824 580 4840 614
rect 4874 580 5853 614
rect 5144 490 5160 524
rect 5194 490 5963 524
rect 5144 266 5160 300
rect 5194 266 5963 300
rect 1360 187 1394 203
rect 0 153 16 187
rect 50 153 1360 187
rect 4824 176 4840 210
rect 4874 176 5853 210
rect 1360 137 1394 153
rect 4426 137 4460 153
rect 7280 103 7857 137
rect 4426 87 4460 103
rect 4504 64 4520 98
rect 4554 64 5963 98
<< viali >>
rect 4760 50462 4794 50496
rect 5080 50350 5114 50384
rect 5720 50260 5754 50294
rect 5720 50036 5754 50070
rect 5080 49946 5114 49980
rect 4680 49834 4714 49868
rect 4600 49672 4634 49706
rect 5080 49560 5114 49594
rect 5720 49470 5754 49504
rect 5720 49246 5754 49280
rect 5080 49156 5114 49190
rect 4520 49044 4554 49078
rect 4760 48882 4794 48916
rect 5000 48770 5034 48804
rect 5720 48680 5754 48714
rect 5720 48456 5754 48490
rect 5000 48366 5034 48400
rect 4680 48254 4714 48288
rect 4600 48092 4634 48126
rect 5000 47980 5034 48014
rect 5720 47890 5754 47924
rect 5720 47666 5754 47700
rect 5000 47576 5034 47610
rect 4520 47464 4554 47498
rect 4760 47302 4794 47336
rect 4920 47190 4954 47224
rect 5720 47100 5754 47134
rect 5720 46876 5754 46910
rect 4920 46786 4954 46820
rect 4680 46674 4714 46708
rect 4600 46512 4634 46546
rect 4920 46400 4954 46434
rect 5720 46310 5754 46344
rect 5720 46086 5754 46120
rect 4920 45996 4954 46030
rect 4520 45884 4554 45918
rect 4760 45722 4794 45756
rect 4840 45610 4874 45644
rect 5720 45520 5754 45554
rect 5720 45296 5754 45330
rect 4840 45206 4874 45240
rect 4680 45094 4714 45128
rect 4600 44932 4634 44966
rect 4840 44820 4874 44854
rect 5720 44730 5754 44764
rect 5720 44506 5754 44540
rect 4840 44416 4874 44450
rect 4520 44304 4554 44338
rect 4760 44142 4794 44176
rect 5080 44030 5114 44064
rect 5640 43940 5674 43974
rect 5640 43716 5674 43750
rect 5080 43626 5114 43660
rect 4680 43514 4714 43548
rect 4600 43352 4634 43386
rect 5080 43240 5114 43274
rect 5640 43150 5674 43184
rect 5640 42926 5674 42960
rect 5080 42836 5114 42870
rect 4520 42724 4554 42758
rect 4760 42562 4794 42596
rect 5000 42450 5034 42484
rect 5640 42360 5674 42394
rect 5640 42136 5674 42170
rect 5000 42046 5034 42080
rect 4680 41934 4714 41968
rect 4600 41772 4634 41806
rect 5000 41660 5034 41694
rect 5640 41570 5674 41604
rect 5640 41346 5674 41380
rect 5000 41256 5034 41290
rect 4520 41144 4554 41178
rect 4760 40982 4794 41016
rect 4920 40870 4954 40904
rect 5640 40780 5674 40814
rect 5640 40556 5674 40590
rect 4920 40466 4954 40500
rect 4680 40354 4714 40388
rect 4600 40192 4634 40226
rect 4920 40080 4954 40114
rect 5640 39990 5674 40024
rect 5640 39766 5674 39800
rect 4920 39676 4954 39710
rect 4520 39564 4554 39598
rect 4760 39402 4794 39436
rect 4840 39290 4874 39324
rect 5640 39200 5674 39234
rect 5640 38976 5674 39010
rect 4840 38886 4874 38920
rect 4680 38774 4714 38808
rect 4600 38612 4634 38646
rect 4840 38500 4874 38534
rect 5640 38410 5674 38444
rect 5640 38186 5674 38220
rect 4840 38096 4874 38130
rect 4520 37984 4554 38018
rect 4760 37822 4794 37856
rect 5080 37710 5114 37744
rect 5560 37620 5594 37654
rect 5560 37396 5594 37430
rect 5080 37306 5114 37340
rect 4680 37194 4714 37228
rect 4600 37032 4634 37066
rect 5080 36920 5114 36954
rect 5560 36830 5594 36864
rect 5560 36606 5594 36640
rect 5080 36516 5114 36550
rect 4520 36404 4554 36438
rect 4760 36242 4794 36276
rect 5000 36130 5034 36164
rect 5560 36040 5594 36074
rect 5560 35816 5594 35850
rect 5000 35726 5034 35760
rect 4680 35614 4714 35648
rect 4600 35452 4634 35486
rect 5000 35340 5034 35374
rect 5560 35250 5594 35284
rect 5560 35026 5594 35060
rect 5000 34936 5034 34970
rect 4520 34824 4554 34858
rect 4760 34662 4794 34696
rect 4920 34550 4954 34584
rect 5560 34460 5594 34494
rect 5560 34236 5594 34270
rect 4920 34146 4954 34180
rect 4680 34034 4714 34068
rect 4600 33872 4634 33906
rect 4920 33760 4954 33794
rect 5560 33670 5594 33704
rect 5560 33446 5594 33480
rect 4920 33356 4954 33390
rect 4520 33244 4554 33278
rect 4760 33082 4794 33116
rect 4840 32970 4874 33004
rect 5560 32880 5594 32914
rect 5560 32656 5594 32690
rect 4840 32566 4874 32600
rect 4680 32454 4714 32488
rect 4600 32292 4634 32326
rect 4840 32180 4874 32214
rect 5560 32090 5594 32124
rect 5560 31866 5594 31900
rect 4840 31776 4874 31810
rect 4520 31664 4554 31698
rect 4760 31502 4794 31536
rect 5080 31390 5114 31424
rect 5480 31300 5514 31334
rect 5480 31076 5514 31110
rect 5080 30986 5114 31020
rect 4680 30874 4714 30908
rect 4600 30712 4634 30746
rect 5080 30600 5114 30634
rect 5480 30510 5514 30544
rect 5480 30286 5514 30320
rect 5080 30196 5114 30230
rect 4520 30084 4554 30118
rect 4760 29922 4794 29956
rect 5000 29810 5034 29844
rect 5480 29720 5514 29754
rect 5480 29496 5514 29530
rect 5000 29406 5034 29440
rect 4680 29294 4714 29328
rect 4600 29132 4634 29166
rect 5000 29020 5034 29054
rect 5480 28930 5514 28964
rect 5480 28706 5514 28740
rect 5000 28616 5034 28650
rect 4520 28504 4554 28538
rect 4760 28342 4794 28376
rect 4920 28230 4954 28264
rect 5480 28140 5514 28174
rect 5480 27916 5514 27950
rect 4920 27826 4954 27860
rect 4680 27714 4714 27748
rect 4600 27552 4634 27586
rect 4920 27440 4954 27474
rect 5480 27350 5514 27384
rect 5480 27126 5514 27160
rect 4920 27036 4954 27070
rect 4520 26924 4554 26958
rect 4760 26762 4794 26796
rect 4840 26650 4874 26684
rect 5480 26560 5514 26594
rect 5480 26336 5514 26370
rect 4840 26246 4874 26280
rect 4680 26134 4714 26168
rect 4600 25972 4634 26006
rect 4840 25860 4874 25894
rect 5480 25770 5514 25804
rect 5480 25546 5514 25580
rect 4840 25456 4874 25490
rect 4520 25344 4554 25378
rect 4760 25182 4794 25216
rect 5080 25070 5114 25104
rect 5400 24980 5434 25014
rect 5400 24756 5434 24790
rect 5080 24666 5114 24700
rect 4680 24554 4714 24588
rect 4600 24392 4634 24426
rect 5080 24280 5114 24314
rect 5400 24190 5434 24224
rect 5400 23966 5434 24000
rect 5080 23876 5114 23910
rect 4520 23764 4554 23798
rect 4760 23602 4794 23636
rect 5000 23490 5034 23524
rect 5400 23400 5434 23434
rect 5400 23176 5434 23210
rect 5000 23086 5034 23120
rect 4680 22974 4714 23008
rect 4600 22812 4634 22846
rect 5000 22700 5034 22734
rect 5400 22610 5434 22644
rect 5400 22386 5434 22420
rect 5000 22296 5034 22330
rect 4520 22184 4554 22218
rect 4760 22022 4794 22056
rect 4920 21910 4954 21944
rect 5400 21820 5434 21854
rect 5400 21596 5434 21630
rect 4920 21506 4954 21540
rect 4680 21394 4714 21428
rect 4600 21232 4634 21266
rect 4920 21120 4954 21154
rect 5400 21030 5434 21064
rect 5400 20806 5434 20840
rect 4920 20716 4954 20750
rect 4520 20604 4554 20638
rect 4760 20442 4794 20476
rect 4840 20330 4874 20364
rect 5400 20240 5434 20274
rect 5400 20016 5434 20050
rect 4840 19926 4874 19960
rect 4680 19814 4714 19848
rect 4600 19652 4634 19686
rect 4840 19540 4874 19574
rect 5400 19450 5434 19484
rect 5400 19226 5434 19260
rect 4840 19136 4874 19170
rect 4520 19024 4554 19058
rect 4760 18862 4794 18896
rect 5080 18750 5114 18784
rect 5320 18660 5354 18694
rect 5320 18436 5354 18470
rect 5080 18346 5114 18380
rect 4680 18234 4714 18268
rect 4600 18072 4634 18106
rect 5080 17960 5114 17994
rect 5320 17870 5354 17904
rect 5320 17646 5354 17680
rect 5080 17556 5114 17590
rect 4520 17444 4554 17478
rect 4760 17282 4794 17316
rect 5000 17170 5034 17204
rect 5320 17080 5354 17114
rect 5320 16856 5354 16890
rect 5000 16766 5034 16800
rect 4680 16654 4714 16688
rect 4600 16492 4634 16526
rect 5000 16380 5034 16414
rect 5320 16290 5354 16324
rect 5320 16066 5354 16100
rect 5000 15976 5034 16010
rect 4520 15864 4554 15898
rect 4760 15702 4794 15736
rect 4920 15590 4954 15624
rect 5320 15500 5354 15534
rect 5320 15276 5354 15310
rect 4920 15186 4954 15220
rect 4680 15074 4714 15108
rect 4600 14912 4634 14946
rect 4920 14800 4954 14834
rect 5320 14710 5354 14744
rect 5320 14486 5354 14520
rect 4920 14396 4954 14430
rect 4520 14284 4554 14318
rect 4760 14122 4794 14156
rect 4840 14010 4874 14044
rect 5320 13920 5354 13954
rect 5320 13696 5354 13730
rect 4840 13606 4874 13640
rect 4680 13494 4714 13528
rect 4600 13332 4634 13366
rect 4840 13220 4874 13254
rect 5320 13130 5354 13164
rect 5320 12906 5354 12940
rect 4840 12816 4874 12850
rect 4520 12704 4554 12738
rect 4760 12542 4794 12576
rect 5080 12430 5114 12464
rect 5240 12340 5274 12374
rect 5240 12116 5274 12150
rect 5080 12026 5114 12060
rect 4680 11914 4714 11948
rect 4600 11752 4634 11786
rect 5080 11640 5114 11674
rect 5240 11550 5274 11584
rect 5240 11326 5274 11360
rect 5080 11236 5114 11270
rect 4520 11124 4554 11158
rect 4760 10962 4794 10996
rect 5000 10850 5034 10884
rect 5240 10760 5274 10794
rect 5240 10536 5274 10570
rect 5000 10446 5034 10480
rect 4680 10334 4714 10368
rect 4600 10172 4634 10206
rect 5000 10060 5034 10094
rect 5240 9970 5274 10004
rect 5240 9746 5274 9780
rect 5000 9656 5034 9690
rect 4520 9544 4554 9578
rect 4760 9382 4794 9416
rect 4920 9270 4954 9304
rect 5240 9180 5274 9214
rect 5240 8956 5274 8990
rect 4920 8866 4954 8900
rect 4680 8754 4714 8788
rect 4600 8592 4634 8626
rect 4920 8480 4954 8514
rect 5240 8390 5274 8424
rect 5240 8166 5274 8200
rect 4920 8076 4954 8110
rect 4520 7964 4554 7998
rect 4760 7802 4794 7836
rect 4426 7763 4460 7797
rect 4840 7690 4874 7724
rect 5240 7600 5274 7634
rect 5240 7376 5274 7410
rect 4840 7286 4874 7320
rect 4426 7213 4460 7247
rect 4680 7174 4714 7208
rect 4600 7012 4634 7046
rect 4426 6973 4460 7007
rect 4840 6900 4874 6934
rect 5240 6810 5274 6844
rect 5240 6586 5274 6620
rect 4840 6496 4874 6530
rect 4426 6423 4460 6457
rect 4520 6384 4554 6418
rect 4760 6222 4794 6256
rect 4426 6183 4460 6217
rect 5080 6110 5114 6144
rect 5160 6020 5194 6054
rect 5160 5796 5194 5830
rect 496 5683 530 5717
rect 844 5683 878 5717
rect 5080 5706 5114 5740
rect 4426 5633 4460 5667
rect 4680 5594 4714 5628
rect 4600 5432 4634 5466
rect 4426 5393 4460 5427
rect 416 5343 450 5377
rect 764 5343 798 5377
rect 5080 5320 5114 5354
rect 5160 5230 5194 5264
rect 5160 5006 5194 5040
rect 336 4893 370 4927
rect 684 4893 718 4927
rect 5080 4916 5114 4950
rect 4426 4843 4460 4877
rect 4520 4804 4554 4838
rect 4760 4642 4794 4676
rect 5000 4530 5034 4564
rect 5160 4440 5194 4474
rect 5160 4216 5194 4250
rect 5000 4126 5034 4160
rect 4680 4014 4714 4048
rect 4600 3852 4634 3886
rect 4426 3813 4460 3847
rect 5000 3740 5034 3774
rect 5160 3650 5194 3684
rect 5160 3426 5194 3460
rect 5000 3336 5034 3370
rect 4426 3263 4460 3297
rect 4520 3224 4554 3258
rect 4760 3062 4794 3096
rect 4426 3023 4460 3057
rect 256 2973 290 3007
rect 1440 2973 1474 3007
rect 4920 2950 4954 2984
rect 5160 2860 5194 2894
rect 5160 2636 5194 2670
rect 176 2523 210 2557
rect 1360 2523 1394 2557
rect 4920 2546 4954 2580
rect 4426 2473 4460 2507
rect 4680 2434 4714 2468
rect 4600 2272 4634 2306
rect 4920 2160 4954 2194
rect 5160 2070 5194 2104
rect 5160 1846 5194 1880
rect 4920 1756 4954 1790
rect 4520 1644 4554 1678
rect 4760 1482 4794 1516
rect 4426 1443 4460 1477
rect 4840 1370 4874 1404
rect 5160 1280 5194 1314
rect 5160 1056 5194 1090
rect 4840 966 4874 1000
rect 4426 893 4460 927
rect 4680 854 4714 888
rect 4600 692 4634 726
rect 4426 653 4460 687
rect 96 603 130 637
rect 1440 603 1474 637
rect 4840 580 4874 614
rect 5160 490 5194 524
rect 5160 266 5194 300
rect 16 153 50 187
rect 1360 153 1394 187
rect 4840 176 4874 210
rect 4426 103 4460 137
rect 4520 64 4554 98
<< metal1 >>
rect 4523 49090 4551 50588
rect 4603 49718 4631 50588
rect 4683 49880 4711 50588
rect 4763 50508 4791 50588
rect 4754 50496 4800 50508
rect 4754 50462 4760 50496
rect 4794 50462 4800 50496
rect 4754 50450 4800 50462
rect 4674 49868 4720 49880
rect 4674 49834 4680 49868
rect 4714 49834 4720 49868
rect 4674 49822 4720 49834
rect 4594 49706 4640 49718
rect 4594 49672 4600 49706
rect 4634 49672 4640 49706
rect 4594 49660 4640 49672
rect 4514 49078 4560 49090
rect 4514 49044 4520 49078
rect 4554 49044 4560 49078
rect 4514 49032 4560 49044
rect 4523 47510 4551 49032
rect 4603 48138 4631 49660
rect 4683 48300 4711 49822
rect 4763 48928 4791 50450
rect 4754 48916 4800 48928
rect 4754 48882 4760 48916
rect 4794 48882 4800 48916
rect 4754 48870 4800 48882
rect 4674 48288 4720 48300
rect 4674 48254 4680 48288
rect 4714 48254 4720 48288
rect 4674 48242 4720 48254
rect 4594 48126 4640 48138
rect 4594 48092 4600 48126
rect 4634 48092 4640 48126
rect 4594 48080 4640 48092
rect 4514 47498 4560 47510
rect 4514 47464 4520 47498
rect 4554 47464 4560 47498
rect 4514 47452 4560 47464
rect 4523 45930 4551 47452
rect 4603 46558 4631 48080
rect 4683 46720 4711 48242
rect 4763 47348 4791 48870
rect 4754 47336 4800 47348
rect 4754 47302 4760 47336
rect 4794 47302 4800 47336
rect 4754 47290 4800 47302
rect 4674 46708 4720 46720
rect 4674 46674 4680 46708
rect 4714 46674 4720 46708
rect 4674 46662 4720 46674
rect 4594 46546 4640 46558
rect 4594 46512 4600 46546
rect 4634 46512 4640 46546
rect 4594 46500 4640 46512
rect 4514 45918 4560 45930
rect 4514 45884 4520 45918
rect 4554 45884 4560 45918
rect 4514 45872 4560 45884
rect 4523 44350 4551 45872
rect 4603 44978 4631 46500
rect 4683 45140 4711 46662
rect 4763 45768 4791 47290
rect 4754 45756 4800 45768
rect 4754 45722 4760 45756
rect 4794 45722 4800 45756
rect 4754 45710 4800 45722
rect 4674 45128 4720 45140
rect 4674 45094 4680 45128
rect 4714 45094 4720 45128
rect 4674 45082 4720 45094
rect 4594 44966 4640 44978
rect 4594 44932 4600 44966
rect 4634 44932 4640 44966
rect 4594 44920 4640 44932
rect 4514 44338 4560 44350
rect 4514 44304 4520 44338
rect 4554 44304 4560 44338
rect 4514 44292 4560 44304
rect 4523 42770 4551 44292
rect 4603 43398 4631 44920
rect 4683 43560 4711 45082
rect 4763 44188 4791 45710
rect 4843 45656 4871 50588
rect 4923 47236 4951 50588
rect 5003 48816 5031 50588
rect 5083 50396 5111 50588
rect 5074 50384 5120 50396
rect 5074 50350 5080 50384
rect 5114 50350 5120 50384
rect 5074 50338 5120 50350
rect 5083 49992 5111 50338
rect 5074 49980 5120 49992
rect 5074 49946 5080 49980
rect 5114 49946 5120 49980
rect 5074 49934 5120 49946
rect 5083 49606 5111 49934
rect 5074 49594 5120 49606
rect 5074 49560 5080 49594
rect 5114 49560 5120 49594
rect 5074 49548 5120 49560
rect 5083 49202 5111 49548
rect 5074 49190 5120 49202
rect 5074 49156 5080 49190
rect 5114 49156 5120 49190
rect 5074 49144 5120 49156
rect 4994 48804 5040 48816
rect 4994 48770 5000 48804
rect 5034 48770 5040 48804
rect 4994 48758 5040 48770
rect 5003 48412 5031 48758
rect 4994 48400 5040 48412
rect 4994 48366 5000 48400
rect 5034 48366 5040 48400
rect 4994 48354 5040 48366
rect 5003 48026 5031 48354
rect 4994 48014 5040 48026
rect 4994 47980 5000 48014
rect 5034 47980 5040 48014
rect 4994 47968 5040 47980
rect 5003 47622 5031 47968
rect 4994 47610 5040 47622
rect 4994 47576 5000 47610
rect 5034 47576 5040 47610
rect 4994 47564 5040 47576
rect 4914 47224 4960 47236
rect 4914 47190 4920 47224
rect 4954 47190 4960 47224
rect 4914 47178 4960 47190
rect 4923 46832 4951 47178
rect 4914 46820 4960 46832
rect 4914 46786 4920 46820
rect 4954 46786 4960 46820
rect 4914 46774 4960 46786
rect 4923 46446 4951 46774
rect 4914 46434 4960 46446
rect 4914 46400 4920 46434
rect 4954 46400 4960 46434
rect 4914 46388 4960 46400
rect 4923 46042 4951 46388
rect 4914 46030 4960 46042
rect 4914 45996 4920 46030
rect 4954 45996 4960 46030
rect 4914 45984 4960 45996
rect 4834 45644 4880 45656
rect 4834 45610 4840 45644
rect 4874 45610 4880 45644
rect 4834 45598 4880 45610
rect 4843 45252 4871 45598
rect 4834 45240 4880 45252
rect 4834 45206 4840 45240
rect 4874 45206 4880 45240
rect 4834 45194 4880 45206
rect 4843 44866 4871 45194
rect 4834 44854 4880 44866
rect 4834 44820 4840 44854
rect 4874 44820 4880 44854
rect 4834 44808 4880 44820
rect 4843 44462 4871 44808
rect 4834 44450 4880 44462
rect 4834 44416 4840 44450
rect 4874 44416 4880 44450
rect 4834 44404 4880 44416
rect 4754 44176 4800 44188
rect 4754 44142 4760 44176
rect 4794 44142 4800 44176
rect 4754 44130 4800 44142
rect 4674 43548 4720 43560
rect 4674 43514 4680 43548
rect 4714 43514 4720 43548
rect 4674 43502 4720 43514
rect 4594 43386 4640 43398
rect 4594 43352 4600 43386
rect 4634 43352 4640 43386
rect 4594 43340 4640 43352
rect 4514 42758 4560 42770
rect 4514 42724 4520 42758
rect 4554 42724 4560 42758
rect 4514 42712 4560 42724
rect 4523 41190 4551 42712
rect 4603 41818 4631 43340
rect 4683 41980 4711 43502
rect 4763 42608 4791 44130
rect 4754 42596 4800 42608
rect 4754 42562 4760 42596
rect 4794 42562 4800 42596
rect 4754 42550 4800 42562
rect 4674 41968 4720 41980
rect 4674 41934 4680 41968
rect 4714 41934 4720 41968
rect 4674 41922 4720 41934
rect 4594 41806 4640 41818
rect 4594 41772 4600 41806
rect 4634 41772 4640 41806
rect 4594 41760 4640 41772
rect 4514 41178 4560 41190
rect 4514 41144 4520 41178
rect 4554 41144 4560 41178
rect 4514 41132 4560 41144
rect 4523 39610 4551 41132
rect 4603 40238 4631 41760
rect 4683 40400 4711 41922
rect 4763 41028 4791 42550
rect 4754 41016 4800 41028
rect 4754 40982 4760 41016
rect 4794 40982 4800 41016
rect 4754 40970 4800 40982
rect 4674 40388 4720 40400
rect 4674 40354 4680 40388
rect 4714 40354 4720 40388
rect 4674 40342 4720 40354
rect 4594 40226 4640 40238
rect 4594 40192 4600 40226
rect 4634 40192 4640 40226
rect 4594 40180 4640 40192
rect 4514 39598 4560 39610
rect 4514 39564 4520 39598
rect 4554 39564 4560 39598
rect 4514 39552 4560 39564
rect 4523 38030 4551 39552
rect 4603 38658 4631 40180
rect 4683 38820 4711 40342
rect 4763 39448 4791 40970
rect 4754 39436 4800 39448
rect 4754 39402 4760 39436
rect 4794 39402 4800 39436
rect 4754 39390 4800 39402
rect 4674 38808 4720 38820
rect 4674 38774 4680 38808
rect 4714 38774 4720 38808
rect 4674 38762 4720 38774
rect 4594 38646 4640 38658
rect 4594 38612 4600 38646
rect 4634 38612 4640 38646
rect 4594 38600 4640 38612
rect 4514 38018 4560 38030
rect 4514 37984 4520 38018
rect 4554 37984 4560 38018
rect 4514 37972 4560 37984
rect 4523 36450 4551 37972
rect 4603 37078 4631 38600
rect 4683 37240 4711 38762
rect 4763 37868 4791 39390
rect 4843 39336 4871 44404
rect 4923 40916 4951 45984
rect 5003 42496 5031 47564
rect 5083 44076 5111 49144
rect 5074 44064 5120 44076
rect 5074 44030 5080 44064
rect 5114 44030 5120 44064
rect 5074 44018 5120 44030
rect 5083 43672 5111 44018
rect 5074 43660 5120 43672
rect 5074 43626 5080 43660
rect 5114 43626 5120 43660
rect 5074 43614 5120 43626
rect 5083 43286 5111 43614
rect 5074 43274 5120 43286
rect 5074 43240 5080 43274
rect 5114 43240 5120 43274
rect 5074 43228 5120 43240
rect 5083 42882 5111 43228
rect 5074 42870 5120 42882
rect 5074 42836 5080 42870
rect 5114 42836 5120 42870
rect 5074 42824 5120 42836
rect 4994 42484 5040 42496
rect 4994 42450 5000 42484
rect 5034 42450 5040 42484
rect 4994 42438 5040 42450
rect 5003 42092 5031 42438
rect 4994 42080 5040 42092
rect 4994 42046 5000 42080
rect 5034 42046 5040 42080
rect 4994 42034 5040 42046
rect 5003 41706 5031 42034
rect 4994 41694 5040 41706
rect 4994 41660 5000 41694
rect 5034 41660 5040 41694
rect 4994 41648 5040 41660
rect 5003 41302 5031 41648
rect 4994 41290 5040 41302
rect 4994 41256 5000 41290
rect 5034 41256 5040 41290
rect 4994 41244 5040 41256
rect 4914 40904 4960 40916
rect 4914 40870 4920 40904
rect 4954 40870 4960 40904
rect 4914 40858 4960 40870
rect 4923 40512 4951 40858
rect 4914 40500 4960 40512
rect 4914 40466 4920 40500
rect 4954 40466 4960 40500
rect 4914 40454 4960 40466
rect 4923 40126 4951 40454
rect 4914 40114 4960 40126
rect 4914 40080 4920 40114
rect 4954 40080 4960 40114
rect 4914 40068 4960 40080
rect 4923 39722 4951 40068
rect 4914 39710 4960 39722
rect 4914 39676 4920 39710
rect 4954 39676 4960 39710
rect 4914 39664 4960 39676
rect 4834 39324 4880 39336
rect 4834 39290 4840 39324
rect 4874 39290 4880 39324
rect 4834 39278 4880 39290
rect 4843 38932 4871 39278
rect 4834 38920 4880 38932
rect 4834 38886 4840 38920
rect 4874 38886 4880 38920
rect 4834 38874 4880 38886
rect 4843 38546 4871 38874
rect 4834 38534 4880 38546
rect 4834 38500 4840 38534
rect 4874 38500 4880 38534
rect 4834 38488 4880 38500
rect 4843 38142 4871 38488
rect 4834 38130 4880 38142
rect 4834 38096 4840 38130
rect 4874 38096 4880 38130
rect 4834 38084 4880 38096
rect 4754 37856 4800 37868
rect 4754 37822 4760 37856
rect 4794 37822 4800 37856
rect 4754 37810 4800 37822
rect 4674 37228 4720 37240
rect 4674 37194 4680 37228
rect 4714 37194 4720 37228
rect 4674 37182 4720 37194
rect 4594 37066 4640 37078
rect 4594 37032 4600 37066
rect 4634 37032 4640 37066
rect 4594 37020 4640 37032
rect 4514 36438 4560 36450
rect 4514 36404 4520 36438
rect 4554 36404 4560 36438
rect 4514 36392 4560 36404
rect 4523 34870 4551 36392
rect 4603 35498 4631 37020
rect 4683 35660 4711 37182
rect 4763 36288 4791 37810
rect 4754 36276 4800 36288
rect 4754 36242 4760 36276
rect 4794 36242 4800 36276
rect 4754 36230 4800 36242
rect 4674 35648 4720 35660
rect 4674 35614 4680 35648
rect 4714 35614 4720 35648
rect 4674 35602 4720 35614
rect 4594 35486 4640 35498
rect 4594 35452 4600 35486
rect 4634 35452 4640 35486
rect 4594 35440 4640 35452
rect 4514 34858 4560 34870
rect 4514 34824 4520 34858
rect 4554 34824 4560 34858
rect 4514 34812 4560 34824
rect 4523 33290 4551 34812
rect 4603 33918 4631 35440
rect 4683 34080 4711 35602
rect 4763 34708 4791 36230
rect 4754 34696 4800 34708
rect 4754 34662 4760 34696
rect 4794 34662 4800 34696
rect 4754 34650 4800 34662
rect 4674 34068 4720 34080
rect 4674 34034 4680 34068
rect 4714 34034 4720 34068
rect 4674 34022 4720 34034
rect 4594 33906 4640 33918
rect 4594 33872 4600 33906
rect 4634 33872 4640 33906
rect 4594 33860 4640 33872
rect 4514 33278 4560 33290
rect 4514 33244 4520 33278
rect 4554 33244 4560 33278
rect 4514 33232 4560 33244
rect 4523 31710 4551 33232
rect 4603 32338 4631 33860
rect 4683 32500 4711 34022
rect 4763 33128 4791 34650
rect 4754 33116 4800 33128
rect 4754 33082 4760 33116
rect 4794 33082 4800 33116
rect 4754 33070 4800 33082
rect 4674 32488 4720 32500
rect 4674 32454 4680 32488
rect 4714 32454 4720 32488
rect 4674 32442 4720 32454
rect 4594 32326 4640 32338
rect 4594 32292 4600 32326
rect 4634 32292 4640 32326
rect 4594 32280 4640 32292
rect 4514 31698 4560 31710
rect 4514 31664 4520 31698
rect 4554 31664 4560 31698
rect 4514 31652 4560 31664
rect 4523 30130 4551 31652
rect 4603 30758 4631 32280
rect 4683 30920 4711 32442
rect 4763 31548 4791 33070
rect 4843 33016 4871 38084
rect 4923 34596 4951 39664
rect 5003 36176 5031 41244
rect 5083 37756 5111 42824
rect 5074 37744 5120 37756
rect 5074 37710 5080 37744
rect 5114 37710 5120 37744
rect 5074 37698 5120 37710
rect 5083 37352 5111 37698
rect 5074 37340 5120 37352
rect 5074 37306 5080 37340
rect 5114 37306 5120 37340
rect 5074 37294 5120 37306
rect 5083 36966 5111 37294
rect 5074 36954 5120 36966
rect 5074 36920 5080 36954
rect 5114 36920 5120 36954
rect 5074 36908 5120 36920
rect 5083 36562 5111 36908
rect 5074 36550 5120 36562
rect 5074 36516 5080 36550
rect 5114 36516 5120 36550
rect 5074 36504 5120 36516
rect 4994 36164 5040 36176
rect 4994 36130 5000 36164
rect 5034 36130 5040 36164
rect 4994 36118 5040 36130
rect 5003 35772 5031 36118
rect 4994 35760 5040 35772
rect 4994 35726 5000 35760
rect 5034 35726 5040 35760
rect 4994 35714 5040 35726
rect 5003 35386 5031 35714
rect 4994 35374 5040 35386
rect 4994 35340 5000 35374
rect 5034 35340 5040 35374
rect 4994 35328 5040 35340
rect 5003 34982 5031 35328
rect 4994 34970 5040 34982
rect 4994 34936 5000 34970
rect 5034 34936 5040 34970
rect 4994 34924 5040 34936
rect 4914 34584 4960 34596
rect 4914 34550 4920 34584
rect 4954 34550 4960 34584
rect 4914 34538 4960 34550
rect 4923 34192 4951 34538
rect 4914 34180 4960 34192
rect 4914 34146 4920 34180
rect 4954 34146 4960 34180
rect 4914 34134 4960 34146
rect 4923 33806 4951 34134
rect 4914 33794 4960 33806
rect 4914 33760 4920 33794
rect 4954 33760 4960 33794
rect 4914 33748 4960 33760
rect 4923 33402 4951 33748
rect 4914 33390 4960 33402
rect 4914 33356 4920 33390
rect 4954 33356 4960 33390
rect 4914 33344 4960 33356
rect 4834 33004 4880 33016
rect 4834 32970 4840 33004
rect 4874 32970 4880 33004
rect 4834 32958 4880 32970
rect 4843 32612 4871 32958
rect 4834 32600 4880 32612
rect 4834 32566 4840 32600
rect 4874 32566 4880 32600
rect 4834 32554 4880 32566
rect 4843 32226 4871 32554
rect 4834 32214 4880 32226
rect 4834 32180 4840 32214
rect 4874 32180 4880 32214
rect 4834 32168 4880 32180
rect 4843 31822 4871 32168
rect 4834 31810 4880 31822
rect 4834 31776 4840 31810
rect 4874 31776 4880 31810
rect 4834 31764 4880 31776
rect 4754 31536 4800 31548
rect 4754 31502 4760 31536
rect 4794 31502 4800 31536
rect 4754 31490 4800 31502
rect 4674 30908 4720 30920
rect 4674 30874 4680 30908
rect 4714 30874 4720 30908
rect 4674 30862 4720 30874
rect 4594 30746 4640 30758
rect 4594 30712 4600 30746
rect 4634 30712 4640 30746
rect 4594 30700 4640 30712
rect 4514 30118 4560 30130
rect 4514 30084 4520 30118
rect 4554 30084 4560 30118
rect 4514 30072 4560 30084
rect 4523 28550 4551 30072
rect 4603 29178 4631 30700
rect 4683 29340 4711 30862
rect 4763 29968 4791 31490
rect 4754 29956 4800 29968
rect 4754 29922 4760 29956
rect 4794 29922 4800 29956
rect 4754 29910 4800 29922
rect 4674 29328 4720 29340
rect 4674 29294 4680 29328
rect 4714 29294 4720 29328
rect 4674 29282 4720 29294
rect 4594 29166 4640 29178
rect 4594 29132 4600 29166
rect 4634 29132 4640 29166
rect 4594 29120 4640 29132
rect 4514 28538 4560 28550
rect 4514 28504 4520 28538
rect 4554 28504 4560 28538
rect 4514 28492 4560 28504
rect 4523 26970 4551 28492
rect 4603 27598 4631 29120
rect 4683 27760 4711 29282
rect 4763 28388 4791 29910
rect 4754 28376 4800 28388
rect 4754 28342 4760 28376
rect 4794 28342 4800 28376
rect 4754 28330 4800 28342
rect 4674 27748 4720 27760
rect 4674 27714 4680 27748
rect 4714 27714 4720 27748
rect 4674 27702 4720 27714
rect 4594 27586 4640 27598
rect 4594 27552 4600 27586
rect 4634 27552 4640 27586
rect 4594 27540 4640 27552
rect 4514 26958 4560 26970
rect 4514 26924 4520 26958
rect 4554 26924 4560 26958
rect 4514 26912 4560 26924
rect 4523 25390 4551 26912
rect 4603 26018 4631 27540
rect 4683 26180 4711 27702
rect 4763 26808 4791 28330
rect 4754 26796 4800 26808
rect 4754 26762 4760 26796
rect 4794 26762 4800 26796
rect 4754 26750 4800 26762
rect 4674 26168 4720 26180
rect 4674 26134 4680 26168
rect 4714 26134 4720 26168
rect 4674 26122 4720 26134
rect 4594 26006 4640 26018
rect 4594 25972 4600 26006
rect 4634 25972 4640 26006
rect 4594 25960 4640 25972
rect 4514 25378 4560 25390
rect 4514 25344 4520 25378
rect 4554 25344 4560 25378
rect 4514 25332 4560 25344
rect 4523 23810 4551 25332
rect 4603 24438 4631 25960
rect 4683 24600 4711 26122
rect 4763 25228 4791 26750
rect 4843 26696 4871 31764
rect 4923 28276 4951 33344
rect 5003 29856 5031 34924
rect 5083 31436 5111 36504
rect 5074 31424 5120 31436
rect 5074 31390 5080 31424
rect 5114 31390 5120 31424
rect 5074 31378 5120 31390
rect 5083 31032 5111 31378
rect 5074 31020 5120 31032
rect 5074 30986 5080 31020
rect 5114 30986 5120 31020
rect 5074 30974 5120 30986
rect 5083 30646 5111 30974
rect 5074 30634 5120 30646
rect 5074 30600 5080 30634
rect 5114 30600 5120 30634
rect 5074 30588 5120 30600
rect 5083 30242 5111 30588
rect 5074 30230 5120 30242
rect 5074 30196 5080 30230
rect 5114 30196 5120 30230
rect 5074 30184 5120 30196
rect 4994 29844 5040 29856
rect 4994 29810 5000 29844
rect 5034 29810 5040 29844
rect 4994 29798 5040 29810
rect 5003 29452 5031 29798
rect 4994 29440 5040 29452
rect 4994 29406 5000 29440
rect 5034 29406 5040 29440
rect 4994 29394 5040 29406
rect 5003 29066 5031 29394
rect 4994 29054 5040 29066
rect 4994 29020 5000 29054
rect 5034 29020 5040 29054
rect 4994 29008 5040 29020
rect 5003 28662 5031 29008
rect 4994 28650 5040 28662
rect 4994 28616 5000 28650
rect 5034 28616 5040 28650
rect 4994 28604 5040 28616
rect 4914 28264 4960 28276
rect 4914 28230 4920 28264
rect 4954 28230 4960 28264
rect 4914 28218 4960 28230
rect 4923 27872 4951 28218
rect 4914 27860 4960 27872
rect 4914 27826 4920 27860
rect 4954 27826 4960 27860
rect 4914 27814 4960 27826
rect 4923 27486 4951 27814
rect 4914 27474 4960 27486
rect 4914 27440 4920 27474
rect 4954 27440 4960 27474
rect 4914 27428 4960 27440
rect 4923 27082 4951 27428
rect 4914 27070 4960 27082
rect 4914 27036 4920 27070
rect 4954 27036 4960 27070
rect 4914 27024 4960 27036
rect 4834 26684 4880 26696
rect 4834 26650 4840 26684
rect 4874 26650 4880 26684
rect 4834 26638 4880 26650
rect 4843 26292 4871 26638
rect 4834 26280 4880 26292
rect 4834 26246 4840 26280
rect 4874 26246 4880 26280
rect 4834 26234 4880 26246
rect 4843 25906 4871 26234
rect 4834 25894 4880 25906
rect 4834 25860 4840 25894
rect 4874 25860 4880 25894
rect 4834 25848 4880 25860
rect 4843 25502 4871 25848
rect 4834 25490 4880 25502
rect 4834 25456 4840 25490
rect 4874 25456 4880 25490
rect 4834 25444 4880 25456
rect 4754 25216 4800 25228
rect 4754 25182 4760 25216
rect 4794 25182 4800 25216
rect 4754 25170 4800 25182
rect 4674 24588 4720 24600
rect 4674 24554 4680 24588
rect 4714 24554 4720 24588
rect 4674 24542 4720 24554
rect 4594 24426 4640 24438
rect 4594 24392 4600 24426
rect 4634 24392 4640 24426
rect 4594 24380 4640 24392
rect 4514 23798 4560 23810
rect 4514 23764 4520 23798
rect 4554 23764 4560 23798
rect 4514 23752 4560 23764
rect 4523 22230 4551 23752
rect 4603 22858 4631 24380
rect 4683 23020 4711 24542
rect 4763 23648 4791 25170
rect 4754 23636 4800 23648
rect 4754 23602 4760 23636
rect 4794 23602 4800 23636
rect 4754 23590 4800 23602
rect 4674 23008 4720 23020
rect 4674 22974 4680 23008
rect 4714 22974 4720 23008
rect 4674 22962 4720 22974
rect 4594 22846 4640 22858
rect 4594 22812 4600 22846
rect 4634 22812 4640 22846
rect 4594 22800 4640 22812
rect 4514 22218 4560 22230
rect 4514 22184 4520 22218
rect 4554 22184 4560 22218
rect 4514 22172 4560 22184
rect 4523 20650 4551 22172
rect 4603 21278 4631 22800
rect 4683 21440 4711 22962
rect 4763 22068 4791 23590
rect 4754 22056 4800 22068
rect 4754 22022 4760 22056
rect 4794 22022 4800 22056
rect 4754 22010 4800 22022
rect 4674 21428 4720 21440
rect 4674 21394 4680 21428
rect 4714 21394 4720 21428
rect 4674 21382 4720 21394
rect 4594 21266 4640 21278
rect 4594 21232 4600 21266
rect 4634 21232 4640 21266
rect 4594 21220 4640 21232
rect 4514 20638 4560 20650
rect 4514 20604 4520 20638
rect 4554 20604 4560 20638
rect 4514 20592 4560 20604
rect 4523 19070 4551 20592
rect 4603 19698 4631 21220
rect 4683 19860 4711 21382
rect 4763 20488 4791 22010
rect 4754 20476 4800 20488
rect 4754 20442 4760 20476
rect 4794 20442 4800 20476
rect 4754 20430 4800 20442
rect 4674 19848 4720 19860
rect 4674 19814 4680 19848
rect 4714 19814 4720 19848
rect 4674 19802 4720 19814
rect 4594 19686 4640 19698
rect 4594 19652 4600 19686
rect 4634 19652 4640 19686
rect 4594 19640 4640 19652
rect 4514 19058 4560 19070
rect 4514 19024 4520 19058
rect 4554 19024 4560 19058
rect 4514 19012 4560 19024
rect 4523 17490 4551 19012
rect 4603 18118 4631 19640
rect 4683 18280 4711 19802
rect 4763 18908 4791 20430
rect 4843 20376 4871 25444
rect 4923 21956 4951 27024
rect 5003 23536 5031 28604
rect 5083 25116 5111 30184
rect 5074 25104 5120 25116
rect 5074 25070 5080 25104
rect 5114 25070 5120 25104
rect 5074 25058 5120 25070
rect 5083 24712 5111 25058
rect 5074 24700 5120 24712
rect 5074 24666 5080 24700
rect 5114 24666 5120 24700
rect 5074 24654 5120 24666
rect 5083 24326 5111 24654
rect 5074 24314 5120 24326
rect 5074 24280 5080 24314
rect 5114 24280 5120 24314
rect 5074 24268 5120 24280
rect 5083 23922 5111 24268
rect 5074 23910 5120 23922
rect 5074 23876 5080 23910
rect 5114 23876 5120 23910
rect 5074 23864 5120 23876
rect 4994 23524 5040 23536
rect 4994 23490 5000 23524
rect 5034 23490 5040 23524
rect 4994 23478 5040 23490
rect 5003 23132 5031 23478
rect 4994 23120 5040 23132
rect 4994 23086 5000 23120
rect 5034 23086 5040 23120
rect 4994 23074 5040 23086
rect 5003 22746 5031 23074
rect 4994 22734 5040 22746
rect 4994 22700 5000 22734
rect 5034 22700 5040 22734
rect 4994 22688 5040 22700
rect 5003 22342 5031 22688
rect 4994 22330 5040 22342
rect 4994 22296 5000 22330
rect 5034 22296 5040 22330
rect 4994 22284 5040 22296
rect 4914 21944 4960 21956
rect 4914 21910 4920 21944
rect 4954 21910 4960 21944
rect 4914 21898 4960 21910
rect 4923 21552 4951 21898
rect 4914 21540 4960 21552
rect 4914 21506 4920 21540
rect 4954 21506 4960 21540
rect 4914 21494 4960 21506
rect 4923 21166 4951 21494
rect 4914 21154 4960 21166
rect 4914 21120 4920 21154
rect 4954 21120 4960 21154
rect 4914 21108 4960 21120
rect 4923 20762 4951 21108
rect 4914 20750 4960 20762
rect 4914 20716 4920 20750
rect 4954 20716 4960 20750
rect 4914 20704 4960 20716
rect 4834 20364 4880 20376
rect 4834 20330 4840 20364
rect 4874 20330 4880 20364
rect 4834 20318 4880 20330
rect 4843 19972 4871 20318
rect 4834 19960 4880 19972
rect 4834 19926 4840 19960
rect 4874 19926 4880 19960
rect 4834 19914 4880 19926
rect 4843 19586 4871 19914
rect 4834 19574 4880 19586
rect 4834 19540 4840 19574
rect 4874 19540 4880 19574
rect 4834 19528 4880 19540
rect 4843 19182 4871 19528
rect 4834 19170 4880 19182
rect 4834 19136 4840 19170
rect 4874 19136 4880 19170
rect 4834 19124 4880 19136
rect 4754 18896 4800 18908
rect 4754 18862 4760 18896
rect 4794 18862 4800 18896
rect 4754 18850 4800 18862
rect 4674 18268 4720 18280
rect 4674 18234 4680 18268
rect 4714 18234 4720 18268
rect 4674 18222 4720 18234
rect 4594 18106 4640 18118
rect 4594 18072 4600 18106
rect 4634 18072 4640 18106
rect 4594 18060 4640 18072
rect 4514 17478 4560 17490
rect 4514 17444 4520 17478
rect 4554 17444 4560 17478
rect 4514 17432 4560 17444
rect 4523 15910 4551 17432
rect 4603 16538 4631 18060
rect 4683 16700 4711 18222
rect 4763 17328 4791 18850
rect 4754 17316 4800 17328
rect 4754 17282 4760 17316
rect 4794 17282 4800 17316
rect 4754 17270 4800 17282
rect 4674 16688 4720 16700
rect 4674 16654 4680 16688
rect 4714 16654 4720 16688
rect 4674 16642 4720 16654
rect 4594 16526 4640 16538
rect 4594 16492 4600 16526
rect 4634 16492 4640 16526
rect 4594 16480 4640 16492
rect 4514 15898 4560 15910
rect 4514 15864 4520 15898
rect 4554 15864 4560 15898
rect 4514 15852 4560 15864
rect 4523 14330 4551 15852
rect 4603 14958 4631 16480
rect 4683 15120 4711 16642
rect 4763 15748 4791 17270
rect 4754 15736 4800 15748
rect 4754 15702 4760 15736
rect 4794 15702 4800 15736
rect 4754 15690 4800 15702
rect 4674 15108 4720 15120
rect 4674 15074 4680 15108
rect 4714 15074 4720 15108
rect 4674 15062 4720 15074
rect 4594 14946 4640 14958
rect 4594 14912 4600 14946
rect 4634 14912 4640 14946
rect 4594 14900 4640 14912
rect 4514 14318 4560 14330
rect 4514 14284 4520 14318
rect 4554 14284 4560 14318
rect 4514 14272 4560 14284
rect 4523 12750 4551 14272
rect 4603 13378 4631 14900
rect 4683 13540 4711 15062
rect 4763 14168 4791 15690
rect 4754 14156 4800 14168
rect 4754 14122 4760 14156
rect 4794 14122 4800 14156
rect 4754 14110 4800 14122
rect 4674 13528 4720 13540
rect 4674 13494 4680 13528
rect 4714 13494 4720 13528
rect 4674 13482 4720 13494
rect 4594 13366 4640 13378
rect 4594 13332 4600 13366
rect 4634 13332 4640 13366
rect 4594 13320 4640 13332
rect 4514 12738 4560 12750
rect 4514 12704 4520 12738
rect 4554 12704 4560 12738
rect 4514 12692 4560 12704
rect 4523 11170 4551 12692
rect 4603 11798 4631 13320
rect 4683 11960 4711 13482
rect 4763 12588 4791 14110
rect 4843 14056 4871 19124
rect 4923 15636 4951 20704
rect 5003 17216 5031 22284
rect 5083 18796 5111 23864
rect 5074 18784 5120 18796
rect 5074 18750 5080 18784
rect 5114 18750 5120 18784
rect 5074 18738 5120 18750
rect 5083 18392 5111 18738
rect 5074 18380 5120 18392
rect 5074 18346 5080 18380
rect 5114 18346 5120 18380
rect 5074 18334 5120 18346
rect 5083 18006 5111 18334
rect 5074 17994 5120 18006
rect 5074 17960 5080 17994
rect 5114 17960 5120 17994
rect 5074 17948 5120 17960
rect 5083 17602 5111 17948
rect 5074 17590 5120 17602
rect 5074 17556 5080 17590
rect 5114 17556 5120 17590
rect 5074 17544 5120 17556
rect 4994 17204 5040 17216
rect 4994 17170 5000 17204
rect 5034 17170 5040 17204
rect 4994 17158 5040 17170
rect 5003 16812 5031 17158
rect 4994 16800 5040 16812
rect 4994 16766 5000 16800
rect 5034 16766 5040 16800
rect 4994 16754 5040 16766
rect 5003 16426 5031 16754
rect 4994 16414 5040 16426
rect 4994 16380 5000 16414
rect 5034 16380 5040 16414
rect 4994 16368 5040 16380
rect 5003 16022 5031 16368
rect 4994 16010 5040 16022
rect 4994 15976 5000 16010
rect 5034 15976 5040 16010
rect 4994 15964 5040 15976
rect 4914 15624 4960 15636
rect 4914 15590 4920 15624
rect 4954 15590 4960 15624
rect 4914 15578 4960 15590
rect 4923 15232 4951 15578
rect 4914 15220 4960 15232
rect 4914 15186 4920 15220
rect 4954 15186 4960 15220
rect 4914 15174 4960 15186
rect 4923 14846 4951 15174
rect 4914 14834 4960 14846
rect 4914 14800 4920 14834
rect 4954 14800 4960 14834
rect 4914 14788 4960 14800
rect 4923 14442 4951 14788
rect 4914 14430 4960 14442
rect 4914 14396 4920 14430
rect 4954 14396 4960 14430
rect 4914 14384 4960 14396
rect 4834 14044 4880 14056
rect 4834 14010 4840 14044
rect 4874 14010 4880 14044
rect 4834 13998 4880 14010
rect 4843 13652 4871 13998
rect 4834 13640 4880 13652
rect 4834 13606 4840 13640
rect 4874 13606 4880 13640
rect 4834 13594 4880 13606
rect 4843 13266 4871 13594
rect 4834 13254 4880 13266
rect 4834 13220 4840 13254
rect 4874 13220 4880 13254
rect 4834 13208 4880 13220
rect 4843 12862 4871 13208
rect 4834 12850 4880 12862
rect 4834 12816 4840 12850
rect 4874 12816 4880 12850
rect 4834 12804 4880 12816
rect 4754 12576 4800 12588
rect 4754 12542 4760 12576
rect 4794 12542 4800 12576
rect 4754 12530 4800 12542
rect 4674 11948 4720 11960
rect 4674 11914 4680 11948
rect 4714 11914 4720 11948
rect 4674 11902 4720 11914
rect 4594 11786 4640 11798
rect 4594 11752 4600 11786
rect 4634 11752 4640 11786
rect 4594 11740 4640 11752
rect 4514 11158 4560 11170
rect 4514 11124 4520 11158
rect 4554 11124 4560 11158
rect 4514 11112 4560 11124
rect 4523 9590 4551 11112
rect 4603 10218 4631 11740
rect 4683 10380 4711 11902
rect 4763 11008 4791 12530
rect 4754 10996 4800 11008
rect 4754 10962 4760 10996
rect 4794 10962 4800 10996
rect 4754 10950 4800 10962
rect 4674 10368 4720 10380
rect 4674 10334 4680 10368
rect 4714 10334 4720 10368
rect 4674 10322 4720 10334
rect 4594 10206 4640 10218
rect 4594 10172 4600 10206
rect 4634 10172 4640 10206
rect 4594 10160 4640 10172
rect 4514 9578 4560 9590
rect 4514 9544 4520 9578
rect 4554 9544 4560 9578
rect 4514 9532 4560 9544
rect 4523 8010 4551 9532
rect 4603 8638 4631 10160
rect 4683 8800 4711 10322
rect 4763 9428 4791 10950
rect 4754 9416 4800 9428
rect 4754 9382 4760 9416
rect 4794 9382 4800 9416
rect 4754 9370 4800 9382
rect 4674 8788 4720 8800
rect 4674 8754 4680 8788
rect 4714 8754 4720 8788
rect 4674 8742 4720 8754
rect 4594 8626 4640 8638
rect 4594 8592 4600 8626
rect 4634 8592 4640 8626
rect 4594 8580 4640 8592
rect 4514 7998 4560 8010
rect 4514 7964 4520 7998
rect 4554 7964 4560 7998
rect 4514 7952 4560 7964
rect 19 199 47 7900
rect 99 649 127 7900
rect 179 2569 207 7900
rect 259 3019 287 7900
rect 339 4939 367 7900
rect 419 5389 447 7900
rect 499 5729 527 7900
rect 4411 7754 4417 7806
rect 4469 7754 4475 7806
rect 4411 7204 4417 7256
rect 4469 7204 4475 7256
rect 4411 6964 4417 7016
rect 4469 6964 4475 7016
rect 4411 6414 4417 6466
rect 4469 6414 4475 6466
rect 4523 6430 4551 7952
rect 4603 7058 4631 8580
rect 4683 7220 4711 8742
rect 4763 7848 4791 9370
rect 4754 7836 4800 7848
rect 4754 7802 4760 7836
rect 4794 7802 4800 7836
rect 4754 7790 4800 7802
rect 4674 7208 4720 7220
rect 4674 7174 4680 7208
rect 4714 7174 4720 7208
rect 4674 7162 4720 7174
rect 4594 7046 4640 7058
rect 4594 7012 4600 7046
rect 4634 7012 4640 7046
rect 4594 7000 4640 7012
rect 4514 6418 4560 6430
rect 4514 6384 4520 6418
rect 4554 6384 4560 6418
rect 4514 6372 4560 6384
rect 4411 6174 4417 6226
rect 4469 6174 4475 6226
rect 490 5717 536 5729
rect 490 5683 496 5717
rect 530 5683 536 5717
rect 490 5671 536 5683
rect 832 5717 890 5723
rect 832 5683 844 5717
rect 878 5683 890 5717
rect 832 5677 890 5683
rect 410 5377 456 5389
rect 410 5343 416 5377
rect 450 5343 456 5377
rect 410 5331 456 5343
rect 330 4927 376 4939
rect 330 4893 336 4927
rect 370 4893 376 4927
rect 330 4881 376 4893
rect 250 3007 296 3019
rect 250 2973 256 3007
rect 290 2973 296 3007
rect 250 2961 296 2973
rect 170 2557 216 2569
rect 170 2523 176 2557
rect 210 2523 216 2557
rect 170 2511 216 2523
rect 90 637 136 649
rect 90 603 96 637
rect 130 603 136 637
rect 90 591 136 603
rect 10 187 56 199
rect 10 153 16 187
rect 50 153 56 187
rect 10 141 56 153
rect 19 0 47 141
rect 99 0 127 591
rect 179 0 207 2511
rect 259 0 287 2961
rect 339 0 367 4881
rect 419 0 447 5331
rect 499 0 527 5671
rect 4411 5624 4417 5676
rect 4469 5624 4475 5676
rect 4411 5384 4417 5436
rect 4469 5384 4475 5436
rect 752 5377 810 5383
rect 752 5343 764 5377
rect 798 5343 810 5377
rect 752 5337 810 5343
rect 672 4927 730 4933
rect 672 4893 684 4927
rect 718 4893 730 4927
rect 672 4887 730 4893
rect 4411 4834 4417 4886
rect 4469 4834 4475 4886
rect 4523 4850 4551 6372
rect 4603 5478 4631 7000
rect 4683 5640 4711 7162
rect 4763 6268 4791 7790
rect 4843 7736 4871 12804
rect 4923 9316 4951 14384
rect 5003 10896 5031 15964
rect 5083 12476 5111 17544
rect 5074 12464 5120 12476
rect 5074 12430 5080 12464
rect 5114 12430 5120 12464
rect 5074 12418 5120 12430
rect 5083 12072 5111 12418
rect 5074 12060 5120 12072
rect 5074 12026 5080 12060
rect 5114 12026 5120 12060
rect 5074 12014 5120 12026
rect 5083 11686 5111 12014
rect 5074 11674 5120 11686
rect 5074 11640 5080 11674
rect 5114 11640 5120 11674
rect 5074 11628 5120 11640
rect 5083 11282 5111 11628
rect 5074 11270 5120 11282
rect 5074 11236 5080 11270
rect 5114 11236 5120 11270
rect 5074 11224 5120 11236
rect 4994 10884 5040 10896
rect 4994 10850 5000 10884
rect 5034 10850 5040 10884
rect 4994 10838 5040 10850
rect 5003 10492 5031 10838
rect 4994 10480 5040 10492
rect 4994 10446 5000 10480
rect 5034 10446 5040 10480
rect 4994 10434 5040 10446
rect 5003 10106 5031 10434
rect 4994 10094 5040 10106
rect 4994 10060 5000 10094
rect 5034 10060 5040 10094
rect 4994 10048 5040 10060
rect 5003 9702 5031 10048
rect 4994 9690 5040 9702
rect 4994 9656 5000 9690
rect 5034 9656 5040 9690
rect 4994 9644 5040 9656
rect 4914 9304 4960 9316
rect 4914 9270 4920 9304
rect 4954 9270 4960 9304
rect 4914 9258 4960 9270
rect 4923 8912 4951 9258
rect 4914 8900 4960 8912
rect 4914 8866 4920 8900
rect 4954 8866 4960 8900
rect 4914 8854 4960 8866
rect 4923 8526 4951 8854
rect 4914 8514 4960 8526
rect 4914 8480 4920 8514
rect 4954 8480 4960 8514
rect 4914 8468 4960 8480
rect 4923 8122 4951 8468
rect 4914 8110 4960 8122
rect 4914 8076 4920 8110
rect 4954 8076 4960 8110
rect 4914 8064 4960 8076
rect 4834 7724 4880 7736
rect 4834 7690 4840 7724
rect 4874 7690 4880 7724
rect 4834 7678 4880 7690
rect 4843 7332 4871 7678
rect 4834 7320 4880 7332
rect 4834 7286 4840 7320
rect 4874 7286 4880 7320
rect 4834 7274 4880 7286
rect 4843 6946 4871 7274
rect 4834 6934 4880 6946
rect 4834 6900 4840 6934
rect 4874 6900 4880 6934
rect 4834 6888 4880 6900
rect 4843 6542 4871 6888
rect 4834 6530 4880 6542
rect 4834 6496 4840 6530
rect 4874 6496 4880 6530
rect 4834 6484 4880 6496
rect 4754 6256 4800 6268
rect 4754 6222 4760 6256
rect 4794 6222 4800 6256
rect 4754 6210 4800 6222
rect 4674 5628 4720 5640
rect 4674 5594 4680 5628
rect 4714 5594 4720 5628
rect 4674 5582 4720 5594
rect 4594 5466 4640 5478
rect 4594 5432 4600 5466
rect 4634 5432 4640 5466
rect 4594 5420 4640 5432
rect 4514 4838 4560 4850
rect 4514 4804 4520 4838
rect 4554 4804 4560 4838
rect 4514 4792 4560 4804
rect 4411 3804 4417 3856
rect 4469 3804 4475 3856
rect 4411 3254 4417 3306
rect 4469 3254 4475 3306
rect 4523 3270 4551 4792
rect 4603 3898 4631 5420
rect 4683 4060 4711 5582
rect 4763 4688 4791 6210
rect 4754 4676 4800 4688
rect 4754 4642 4760 4676
rect 4794 4642 4800 4676
rect 4754 4630 4800 4642
rect 4674 4048 4720 4060
rect 4674 4014 4680 4048
rect 4714 4014 4720 4048
rect 4674 4002 4720 4014
rect 4594 3886 4640 3898
rect 4594 3852 4600 3886
rect 4634 3852 4640 3886
rect 4594 3840 4640 3852
rect 4514 3258 4560 3270
rect 4514 3224 4520 3258
rect 4554 3224 4560 3258
rect 4514 3212 4560 3224
rect 4411 3014 4417 3066
rect 4469 3014 4475 3066
rect 1428 3007 1486 3013
rect 1428 2973 1440 3007
rect 1474 2973 1486 3007
rect 1428 2967 1486 2973
rect 1348 2557 1406 2563
rect 1348 2523 1360 2557
rect 1394 2523 1406 2557
rect 1348 2517 1406 2523
rect 4411 2464 4417 2516
rect 4469 2464 4475 2516
rect 4523 1690 4551 3212
rect 4603 2318 4631 3840
rect 4683 2480 4711 4002
rect 4763 3108 4791 4630
rect 4754 3096 4800 3108
rect 4754 3062 4760 3096
rect 4794 3062 4800 3096
rect 4754 3050 4800 3062
rect 4674 2468 4720 2480
rect 4674 2434 4680 2468
rect 4714 2434 4720 2468
rect 4674 2422 4720 2434
rect 4594 2306 4640 2318
rect 4594 2272 4600 2306
rect 4634 2272 4640 2306
rect 4594 2260 4640 2272
rect 4514 1678 4560 1690
rect 4514 1644 4520 1678
rect 4554 1644 4560 1678
rect 4514 1632 4560 1644
rect 4411 1434 4417 1486
rect 4469 1434 4475 1486
rect 4411 884 4417 936
rect 4469 884 4475 936
rect 4411 644 4417 696
rect 4469 644 4475 696
rect 1428 637 1486 643
rect 1428 603 1440 637
rect 1474 603 1486 637
rect 1428 597 1486 603
rect 4523 198 4551 1632
rect 4603 738 4631 2260
rect 4683 988 4711 2422
rect 4763 1528 4791 3050
rect 4843 2568 4871 6484
rect 4923 2996 4951 8064
rect 5003 4576 5031 9644
rect 5083 6156 5111 11224
rect 5074 6144 5120 6156
rect 5074 6110 5080 6144
rect 5114 6110 5120 6144
rect 5074 6098 5120 6110
rect 5083 5752 5111 6098
rect 5163 6066 5191 50588
rect 5243 12386 5271 50588
rect 5323 18706 5351 50588
rect 5403 25026 5431 50588
rect 5483 31346 5511 50588
rect 5563 37666 5591 50588
rect 5643 43986 5671 50588
rect 5723 50306 5751 50588
rect 5714 50294 5760 50306
rect 5714 50260 5720 50294
rect 5754 50260 5760 50294
rect 5714 50248 5760 50260
rect 5723 50082 5751 50248
rect 6051 50214 6097 50516
rect 6475 50214 6523 50574
rect 6907 50214 6955 50574
rect 6042 50162 6048 50214
rect 6100 50162 6106 50214
rect 6467 50162 6473 50214
rect 6525 50162 6531 50214
rect 6899 50162 6905 50214
rect 6957 50162 6963 50214
rect 7299 50191 7327 50560
rect 7695 50191 7723 50560
rect 5714 50070 5760 50082
rect 5714 50036 5720 50070
rect 5754 50036 5760 50070
rect 5714 50024 5760 50036
rect 5723 49516 5751 50024
rect 6051 49840 6097 50162
rect 6042 49788 6048 49840
rect 6100 49788 6106 49840
rect 5714 49504 5760 49516
rect 5714 49470 5720 49504
rect 5754 49470 5760 49504
rect 5714 49458 5760 49470
rect 5723 49292 5751 49458
rect 6051 49424 6097 49788
rect 6475 49782 6523 50162
rect 6907 49782 6955 50162
rect 7281 50139 7287 50191
rect 7339 50139 7345 50191
rect 7677 50139 7683 50191
rect 7735 50139 7741 50191
rect 7299 49796 7327 50139
rect 7695 49796 7723 50139
rect 6467 49730 6473 49782
rect 6525 49730 6531 49782
rect 6899 49730 6905 49782
rect 6957 49730 6963 49782
rect 7281 49744 7287 49796
rect 7339 49744 7345 49796
rect 7677 49744 7683 49796
rect 7735 49744 7741 49796
rect 6475 49424 6523 49730
rect 6907 49424 6955 49730
rect 6042 49372 6048 49424
rect 6100 49372 6106 49424
rect 6467 49372 6473 49424
rect 6525 49372 6531 49424
rect 6899 49372 6905 49424
rect 6957 49372 6963 49424
rect 7299 49401 7327 49744
rect 7695 49401 7723 49744
rect 5714 49280 5760 49292
rect 5714 49246 5720 49280
rect 5754 49246 5760 49280
rect 5714 49234 5760 49246
rect 5723 48726 5751 49234
rect 6051 49050 6097 49372
rect 6042 48998 6048 49050
rect 6100 48998 6106 49050
rect 5714 48714 5760 48726
rect 5714 48680 5720 48714
rect 5754 48680 5760 48714
rect 5714 48668 5760 48680
rect 5723 48502 5751 48668
rect 6051 48634 6097 48998
rect 6475 48992 6523 49372
rect 6907 48992 6955 49372
rect 7281 49349 7287 49401
rect 7339 49349 7345 49401
rect 7677 49349 7683 49401
rect 7735 49349 7741 49401
rect 7299 49006 7327 49349
rect 7695 49006 7723 49349
rect 6467 48940 6473 48992
rect 6525 48940 6531 48992
rect 6899 48940 6905 48992
rect 6957 48940 6963 48992
rect 7281 48954 7287 49006
rect 7339 48954 7345 49006
rect 7677 48954 7683 49006
rect 7735 48954 7741 49006
rect 6475 48634 6523 48940
rect 6907 48634 6955 48940
rect 6042 48582 6048 48634
rect 6100 48582 6106 48634
rect 6467 48582 6473 48634
rect 6525 48582 6531 48634
rect 6899 48582 6905 48634
rect 6957 48582 6963 48634
rect 7299 48611 7327 48954
rect 7695 48611 7723 48954
rect 5714 48490 5760 48502
rect 5714 48456 5720 48490
rect 5754 48456 5760 48490
rect 5714 48444 5760 48456
rect 5723 47936 5751 48444
rect 6051 48260 6097 48582
rect 6042 48208 6048 48260
rect 6100 48208 6106 48260
rect 5714 47924 5760 47936
rect 5714 47890 5720 47924
rect 5754 47890 5760 47924
rect 5714 47878 5760 47890
rect 5723 47712 5751 47878
rect 6051 47844 6097 48208
rect 6475 48202 6523 48582
rect 6907 48202 6955 48582
rect 7281 48559 7287 48611
rect 7339 48559 7345 48611
rect 7677 48559 7683 48611
rect 7735 48559 7741 48611
rect 7299 48216 7327 48559
rect 7695 48216 7723 48559
rect 6467 48150 6473 48202
rect 6525 48150 6531 48202
rect 6899 48150 6905 48202
rect 6957 48150 6963 48202
rect 7281 48164 7287 48216
rect 7339 48164 7345 48216
rect 7677 48164 7683 48216
rect 7735 48164 7741 48216
rect 6475 47844 6523 48150
rect 6907 47844 6955 48150
rect 6042 47792 6048 47844
rect 6100 47792 6106 47844
rect 6467 47792 6473 47844
rect 6525 47792 6531 47844
rect 6899 47792 6905 47844
rect 6957 47792 6963 47844
rect 7299 47821 7327 48164
rect 7695 47821 7723 48164
rect 5714 47700 5760 47712
rect 5714 47666 5720 47700
rect 5754 47666 5760 47700
rect 5714 47654 5760 47666
rect 5723 47146 5751 47654
rect 6051 47470 6097 47792
rect 6042 47418 6048 47470
rect 6100 47418 6106 47470
rect 5714 47134 5760 47146
rect 5714 47100 5720 47134
rect 5754 47100 5760 47134
rect 5714 47088 5760 47100
rect 5723 46922 5751 47088
rect 6051 47054 6097 47418
rect 6475 47412 6523 47792
rect 6907 47412 6955 47792
rect 7281 47769 7287 47821
rect 7339 47769 7345 47821
rect 7677 47769 7683 47821
rect 7735 47769 7741 47821
rect 7299 47426 7327 47769
rect 7695 47426 7723 47769
rect 6467 47360 6473 47412
rect 6525 47360 6531 47412
rect 6899 47360 6905 47412
rect 6957 47360 6963 47412
rect 7281 47374 7287 47426
rect 7339 47374 7345 47426
rect 7677 47374 7683 47426
rect 7735 47374 7741 47426
rect 6475 47054 6523 47360
rect 6907 47054 6955 47360
rect 6042 47002 6048 47054
rect 6100 47002 6106 47054
rect 6467 47002 6473 47054
rect 6525 47002 6531 47054
rect 6899 47002 6905 47054
rect 6957 47002 6963 47054
rect 7299 47031 7327 47374
rect 7695 47031 7723 47374
rect 5714 46910 5760 46922
rect 5714 46876 5720 46910
rect 5754 46876 5760 46910
rect 5714 46864 5760 46876
rect 5723 46356 5751 46864
rect 6051 46680 6097 47002
rect 6042 46628 6048 46680
rect 6100 46628 6106 46680
rect 5714 46344 5760 46356
rect 5714 46310 5720 46344
rect 5754 46310 5760 46344
rect 5714 46298 5760 46310
rect 5723 46132 5751 46298
rect 6051 46264 6097 46628
rect 6475 46622 6523 47002
rect 6907 46622 6955 47002
rect 7281 46979 7287 47031
rect 7339 46979 7345 47031
rect 7677 46979 7683 47031
rect 7735 46979 7741 47031
rect 7299 46636 7327 46979
rect 7695 46636 7723 46979
rect 6467 46570 6473 46622
rect 6525 46570 6531 46622
rect 6899 46570 6905 46622
rect 6957 46570 6963 46622
rect 7281 46584 7287 46636
rect 7339 46584 7345 46636
rect 7677 46584 7683 46636
rect 7735 46584 7741 46636
rect 6475 46264 6523 46570
rect 6907 46264 6955 46570
rect 6042 46212 6048 46264
rect 6100 46212 6106 46264
rect 6467 46212 6473 46264
rect 6525 46212 6531 46264
rect 6899 46212 6905 46264
rect 6957 46212 6963 46264
rect 7299 46241 7327 46584
rect 7695 46241 7723 46584
rect 5714 46120 5760 46132
rect 5714 46086 5720 46120
rect 5754 46086 5760 46120
rect 5714 46074 5760 46086
rect 5723 45566 5751 46074
rect 6051 45890 6097 46212
rect 6042 45838 6048 45890
rect 6100 45838 6106 45890
rect 5714 45554 5760 45566
rect 5714 45520 5720 45554
rect 5754 45520 5760 45554
rect 5714 45508 5760 45520
rect 5723 45342 5751 45508
rect 6051 45474 6097 45838
rect 6475 45832 6523 46212
rect 6907 45832 6955 46212
rect 7281 46189 7287 46241
rect 7339 46189 7345 46241
rect 7677 46189 7683 46241
rect 7735 46189 7741 46241
rect 7299 45846 7327 46189
rect 7695 45846 7723 46189
rect 6467 45780 6473 45832
rect 6525 45780 6531 45832
rect 6899 45780 6905 45832
rect 6957 45780 6963 45832
rect 7281 45794 7287 45846
rect 7339 45794 7345 45846
rect 7677 45794 7683 45846
rect 7735 45794 7741 45846
rect 6475 45474 6523 45780
rect 6907 45474 6955 45780
rect 6042 45422 6048 45474
rect 6100 45422 6106 45474
rect 6467 45422 6473 45474
rect 6525 45422 6531 45474
rect 6899 45422 6905 45474
rect 6957 45422 6963 45474
rect 7299 45451 7327 45794
rect 7695 45451 7723 45794
rect 5714 45330 5760 45342
rect 5714 45296 5720 45330
rect 5754 45296 5760 45330
rect 5714 45284 5760 45296
rect 5723 44776 5751 45284
rect 6051 45100 6097 45422
rect 6042 45048 6048 45100
rect 6100 45048 6106 45100
rect 5714 44764 5760 44776
rect 5714 44730 5720 44764
rect 5754 44730 5760 44764
rect 5714 44718 5760 44730
rect 5723 44552 5751 44718
rect 6051 44684 6097 45048
rect 6475 45042 6523 45422
rect 6907 45042 6955 45422
rect 7281 45399 7287 45451
rect 7339 45399 7345 45451
rect 7677 45399 7683 45451
rect 7735 45399 7741 45451
rect 7299 45056 7327 45399
rect 7695 45056 7723 45399
rect 6467 44990 6473 45042
rect 6525 44990 6531 45042
rect 6899 44990 6905 45042
rect 6957 44990 6963 45042
rect 7281 45004 7287 45056
rect 7339 45004 7345 45056
rect 7677 45004 7683 45056
rect 7735 45004 7741 45056
rect 6475 44684 6523 44990
rect 6907 44684 6955 44990
rect 6042 44632 6048 44684
rect 6100 44632 6106 44684
rect 6467 44632 6473 44684
rect 6525 44632 6531 44684
rect 6899 44632 6905 44684
rect 6957 44632 6963 44684
rect 7299 44661 7327 45004
rect 7695 44661 7723 45004
rect 5714 44540 5760 44552
rect 5714 44506 5720 44540
rect 5754 44506 5760 44540
rect 5714 44494 5760 44506
rect 5634 43974 5680 43986
rect 5634 43940 5640 43974
rect 5674 43940 5680 43974
rect 5634 43928 5680 43940
rect 5643 43762 5671 43928
rect 5634 43750 5680 43762
rect 5634 43716 5640 43750
rect 5674 43716 5680 43750
rect 5634 43704 5680 43716
rect 5643 43196 5671 43704
rect 5634 43184 5680 43196
rect 5634 43150 5640 43184
rect 5674 43150 5680 43184
rect 5634 43138 5680 43150
rect 5643 42972 5671 43138
rect 5634 42960 5680 42972
rect 5634 42926 5640 42960
rect 5674 42926 5680 42960
rect 5634 42914 5680 42926
rect 5643 42406 5671 42914
rect 5634 42394 5680 42406
rect 5634 42360 5640 42394
rect 5674 42360 5680 42394
rect 5634 42348 5680 42360
rect 5643 42182 5671 42348
rect 5634 42170 5680 42182
rect 5634 42136 5640 42170
rect 5674 42136 5680 42170
rect 5634 42124 5680 42136
rect 5643 41616 5671 42124
rect 5634 41604 5680 41616
rect 5634 41570 5640 41604
rect 5674 41570 5680 41604
rect 5634 41558 5680 41570
rect 5643 41392 5671 41558
rect 5634 41380 5680 41392
rect 5634 41346 5640 41380
rect 5674 41346 5680 41380
rect 5634 41334 5680 41346
rect 5643 40826 5671 41334
rect 5634 40814 5680 40826
rect 5634 40780 5640 40814
rect 5674 40780 5680 40814
rect 5634 40768 5680 40780
rect 5643 40602 5671 40768
rect 5634 40590 5680 40602
rect 5634 40556 5640 40590
rect 5674 40556 5680 40590
rect 5634 40544 5680 40556
rect 5643 40036 5671 40544
rect 5634 40024 5680 40036
rect 5634 39990 5640 40024
rect 5674 39990 5680 40024
rect 5634 39978 5680 39990
rect 5643 39812 5671 39978
rect 5634 39800 5680 39812
rect 5634 39766 5640 39800
rect 5674 39766 5680 39800
rect 5634 39754 5680 39766
rect 5643 39246 5671 39754
rect 5634 39234 5680 39246
rect 5634 39200 5640 39234
rect 5674 39200 5680 39234
rect 5634 39188 5680 39200
rect 5643 39022 5671 39188
rect 5634 39010 5680 39022
rect 5634 38976 5640 39010
rect 5674 38976 5680 39010
rect 5634 38964 5680 38976
rect 5643 38456 5671 38964
rect 5634 38444 5680 38456
rect 5634 38410 5640 38444
rect 5674 38410 5680 38444
rect 5634 38398 5680 38410
rect 5643 38232 5671 38398
rect 5634 38220 5680 38232
rect 5634 38186 5640 38220
rect 5674 38186 5680 38220
rect 5634 38174 5680 38186
rect 5554 37654 5600 37666
rect 5554 37620 5560 37654
rect 5594 37620 5600 37654
rect 5554 37608 5600 37620
rect 5563 37442 5591 37608
rect 5554 37430 5600 37442
rect 5554 37396 5560 37430
rect 5594 37396 5600 37430
rect 5554 37384 5600 37396
rect 5563 36876 5591 37384
rect 5554 36864 5600 36876
rect 5554 36830 5560 36864
rect 5594 36830 5600 36864
rect 5554 36818 5600 36830
rect 5563 36652 5591 36818
rect 5554 36640 5600 36652
rect 5554 36606 5560 36640
rect 5594 36606 5600 36640
rect 5554 36594 5600 36606
rect 5563 36086 5591 36594
rect 5554 36074 5600 36086
rect 5554 36040 5560 36074
rect 5594 36040 5600 36074
rect 5554 36028 5600 36040
rect 5563 35862 5591 36028
rect 5554 35850 5600 35862
rect 5554 35816 5560 35850
rect 5594 35816 5600 35850
rect 5554 35804 5600 35816
rect 5563 35296 5591 35804
rect 5554 35284 5600 35296
rect 5554 35250 5560 35284
rect 5594 35250 5600 35284
rect 5554 35238 5600 35250
rect 5563 35072 5591 35238
rect 5554 35060 5600 35072
rect 5554 35026 5560 35060
rect 5594 35026 5600 35060
rect 5554 35014 5600 35026
rect 5563 34506 5591 35014
rect 5554 34494 5600 34506
rect 5554 34460 5560 34494
rect 5594 34460 5600 34494
rect 5554 34448 5600 34460
rect 5563 34282 5591 34448
rect 5554 34270 5600 34282
rect 5554 34236 5560 34270
rect 5594 34236 5600 34270
rect 5554 34224 5600 34236
rect 5563 33716 5591 34224
rect 5554 33704 5600 33716
rect 5554 33670 5560 33704
rect 5594 33670 5600 33704
rect 5554 33658 5600 33670
rect 5563 33492 5591 33658
rect 5554 33480 5600 33492
rect 5554 33446 5560 33480
rect 5594 33446 5600 33480
rect 5554 33434 5600 33446
rect 5563 32926 5591 33434
rect 5554 32914 5600 32926
rect 5554 32880 5560 32914
rect 5594 32880 5600 32914
rect 5554 32868 5600 32880
rect 5563 32702 5591 32868
rect 5554 32690 5600 32702
rect 5554 32656 5560 32690
rect 5594 32656 5600 32690
rect 5554 32644 5600 32656
rect 5563 32136 5591 32644
rect 5554 32124 5600 32136
rect 5554 32090 5560 32124
rect 5594 32090 5600 32124
rect 5554 32078 5600 32090
rect 5563 31912 5591 32078
rect 5554 31900 5600 31912
rect 5554 31866 5560 31900
rect 5594 31866 5600 31900
rect 5554 31854 5600 31866
rect 5474 31334 5520 31346
rect 5474 31300 5480 31334
rect 5514 31300 5520 31334
rect 5474 31288 5520 31300
rect 5483 31122 5511 31288
rect 5474 31110 5520 31122
rect 5474 31076 5480 31110
rect 5514 31076 5520 31110
rect 5474 31064 5520 31076
rect 5483 30556 5511 31064
rect 5474 30544 5520 30556
rect 5474 30510 5480 30544
rect 5514 30510 5520 30544
rect 5474 30498 5520 30510
rect 5483 30332 5511 30498
rect 5474 30320 5520 30332
rect 5474 30286 5480 30320
rect 5514 30286 5520 30320
rect 5474 30274 5520 30286
rect 5483 29766 5511 30274
rect 5474 29754 5520 29766
rect 5474 29720 5480 29754
rect 5514 29720 5520 29754
rect 5474 29708 5520 29720
rect 5483 29542 5511 29708
rect 5474 29530 5520 29542
rect 5474 29496 5480 29530
rect 5514 29496 5520 29530
rect 5474 29484 5520 29496
rect 5483 28976 5511 29484
rect 5474 28964 5520 28976
rect 5474 28930 5480 28964
rect 5514 28930 5520 28964
rect 5474 28918 5520 28930
rect 5483 28752 5511 28918
rect 5474 28740 5520 28752
rect 5474 28706 5480 28740
rect 5514 28706 5520 28740
rect 5474 28694 5520 28706
rect 5483 28186 5511 28694
rect 5474 28174 5520 28186
rect 5474 28140 5480 28174
rect 5514 28140 5520 28174
rect 5474 28128 5520 28140
rect 5483 27962 5511 28128
rect 5474 27950 5520 27962
rect 5474 27916 5480 27950
rect 5514 27916 5520 27950
rect 5474 27904 5520 27916
rect 5483 27396 5511 27904
rect 5474 27384 5520 27396
rect 5474 27350 5480 27384
rect 5514 27350 5520 27384
rect 5474 27338 5520 27350
rect 5483 27172 5511 27338
rect 5474 27160 5520 27172
rect 5474 27126 5480 27160
rect 5514 27126 5520 27160
rect 5474 27114 5520 27126
rect 5483 26606 5511 27114
rect 5474 26594 5520 26606
rect 5474 26560 5480 26594
rect 5514 26560 5520 26594
rect 5474 26548 5520 26560
rect 5483 26382 5511 26548
rect 5474 26370 5520 26382
rect 5474 26336 5480 26370
rect 5514 26336 5520 26370
rect 5474 26324 5520 26336
rect 5483 25816 5511 26324
rect 5474 25804 5520 25816
rect 5474 25770 5480 25804
rect 5514 25770 5520 25804
rect 5474 25758 5520 25770
rect 5483 25592 5511 25758
rect 5474 25580 5520 25592
rect 5474 25546 5480 25580
rect 5514 25546 5520 25580
rect 5474 25534 5520 25546
rect 5394 25014 5440 25026
rect 5394 24980 5400 25014
rect 5434 24980 5440 25014
rect 5394 24968 5440 24980
rect 5403 24802 5431 24968
rect 5394 24790 5440 24802
rect 5394 24756 5400 24790
rect 5434 24756 5440 24790
rect 5394 24744 5440 24756
rect 5403 24236 5431 24744
rect 5394 24224 5440 24236
rect 5394 24190 5400 24224
rect 5434 24190 5440 24224
rect 5394 24178 5440 24190
rect 5403 24012 5431 24178
rect 5394 24000 5440 24012
rect 5394 23966 5400 24000
rect 5434 23966 5440 24000
rect 5394 23954 5440 23966
rect 5403 23446 5431 23954
rect 5394 23434 5440 23446
rect 5394 23400 5400 23434
rect 5434 23400 5440 23434
rect 5394 23388 5440 23400
rect 5403 23222 5431 23388
rect 5394 23210 5440 23222
rect 5394 23176 5400 23210
rect 5434 23176 5440 23210
rect 5394 23164 5440 23176
rect 5403 22656 5431 23164
rect 5394 22644 5440 22656
rect 5394 22610 5400 22644
rect 5434 22610 5440 22644
rect 5394 22598 5440 22610
rect 5403 22432 5431 22598
rect 5394 22420 5440 22432
rect 5394 22386 5400 22420
rect 5434 22386 5440 22420
rect 5394 22374 5440 22386
rect 5403 21866 5431 22374
rect 5394 21854 5440 21866
rect 5394 21820 5400 21854
rect 5434 21820 5440 21854
rect 5394 21808 5440 21820
rect 5403 21642 5431 21808
rect 5394 21630 5440 21642
rect 5394 21596 5400 21630
rect 5434 21596 5440 21630
rect 5394 21584 5440 21596
rect 5403 21076 5431 21584
rect 5394 21064 5440 21076
rect 5394 21030 5400 21064
rect 5434 21030 5440 21064
rect 5394 21018 5440 21030
rect 5403 20852 5431 21018
rect 5394 20840 5440 20852
rect 5394 20806 5400 20840
rect 5434 20806 5440 20840
rect 5394 20794 5440 20806
rect 5403 20286 5431 20794
rect 5394 20274 5440 20286
rect 5394 20240 5400 20274
rect 5434 20240 5440 20274
rect 5394 20228 5440 20240
rect 5403 20062 5431 20228
rect 5394 20050 5440 20062
rect 5394 20016 5400 20050
rect 5434 20016 5440 20050
rect 5394 20004 5440 20016
rect 5403 19496 5431 20004
rect 5394 19484 5440 19496
rect 5394 19450 5400 19484
rect 5434 19450 5440 19484
rect 5394 19438 5440 19450
rect 5403 19272 5431 19438
rect 5394 19260 5440 19272
rect 5394 19226 5400 19260
rect 5434 19226 5440 19260
rect 5394 19214 5440 19226
rect 5314 18694 5360 18706
rect 5314 18660 5320 18694
rect 5354 18660 5360 18694
rect 5314 18648 5360 18660
rect 5323 18482 5351 18648
rect 5314 18470 5360 18482
rect 5314 18436 5320 18470
rect 5354 18436 5360 18470
rect 5314 18424 5360 18436
rect 5323 17916 5351 18424
rect 5314 17904 5360 17916
rect 5314 17870 5320 17904
rect 5354 17870 5360 17904
rect 5314 17858 5360 17870
rect 5323 17692 5351 17858
rect 5314 17680 5360 17692
rect 5314 17646 5320 17680
rect 5354 17646 5360 17680
rect 5314 17634 5360 17646
rect 5323 17126 5351 17634
rect 5314 17114 5360 17126
rect 5314 17080 5320 17114
rect 5354 17080 5360 17114
rect 5314 17068 5360 17080
rect 5323 16902 5351 17068
rect 5314 16890 5360 16902
rect 5314 16856 5320 16890
rect 5354 16856 5360 16890
rect 5314 16844 5360 16856
rect 5323 16336 5351 16844
rect 5314 16324 5360 16336
rect 5314 16290 5320 16324
rect 5354 16290 5360 16324
rect 5314 16278 5360 16290
rect 5323 16112 5351 16278
rect 5314 16100 5360 16112
rect 5314 16066 5320 16100
rect 5354 16066 5360 16100
rect 5314 16054 5360 16066
rect 5323 15546 5351 16054
rect 5314 15534 5360 15546
rect 5314 15500 5320 15534
rect 5354 15500 5360 15534
rect 5314 15488 5360 15500
rect 5323 15322 5351 15488
rect 5314 15310 5360 15322
rect 5314 15276 5320 15310
rect 5354 15276 5360 15310
rect 5314 15264 5360 15276
rect 5323 14756 5351 15264
rect 5314 14744 5360 14756
rect 5314 14710 5320 14744
rect 5354 14710 5360 14744
rect 5314 14698 5360 14710
rect 5323 14532 5351 14698
rect 5314 14520 5360 14532
rect 5314 14486 5320 14520
rect 5354 14486 5360 14520
rect 5314 14474 5360 14486
rect 5323 13966 5351 14474
rect 5314 13954 5360 13966
rect 5314 13920 5320 13954
rect 5354 13920 5360 13954
rect 5314 13908 5360 13920
rect 5323 13742 5351 13908
rect 5314 13730 5360 13742
rect 5314 13696 5320 13730
rect 5354 13696 5360 13730
rect 5314 13684 5360 13696
rect 5323 13176 5351 13684
rect 5314 13164 5360 13176
rect 5314 13130 5320 13164
rect 5354 13130 5360 13164
rect 5314 13118 5360 13130
rect 5323 12952 5351 13118
rect 5314 12940 5360 12952
rect 5314 12906 5320 12940
rect 5354 12906 5360 12940
rect 5314 12894 5360 12906
rect 5234 12374 5280 12386
rect 5234 12340 5240 12374
rect 5274 12340 5280 12374
rect 5234 12328 5280 12340
rect 5243 12162 5271 12328
rect 5234 12150 5280 12162
rect 5234 12116 5240 12150
rect 5274 12116 5280 12150
rect 5234 12104 5280 12116
rect 5243 11596 5271 12104
rect 5234 11584 5280 11596
rect 5234 11550 5240 11584
rect 5274 11550 5280 11584
rect 5234 11538 5280 11550
rect 5243 11372 5271 11538
rect 5234 11360 5280 11372
rect 5234 11326 5240 11360
rect 5274 11326 5280 11360
rect 5234 11314 5280 11326
rect 5243 10806 5271 11314
rect 5234 10794 5280 10806
rect 5234 10760 5240 10794
rect 5274 10760 5280 10794
rect 5234 10748 5280 10760
rect 5243 10582 5271 10748
rect 5234 10570 5280 10582
rect 5234 10536 5240 10570
rect 5274 10536 5280 10570
rect 5234 10524 5280 10536
rect 5243 10016 5271 10524
rect 5234 10004 5280 10016
rect 5234 9970 5240 10004
rect 5274 9970 5280 10004
rect 5234 9958 5280 9970
rect 5243 9792 5271 9958
rect 5234 9780 5280 9792
rect 5234 9746 5240 9780
rect 5274 9746 5280 9780
rect 5234 9734 5280 9746
rect 5243 9226 5271 9734
rect 5234 9214 5280 9226
rect 5234 9180 5240 9214
rect 5274 9180 5280 9214
rect 5234 9168 5280 9180
rect 5243 9002 5271 9168
rect 5234 8990 5280 9002
rect 5234 8956 5240 8990
rect 5274 8956 5280 8990
rect 5234 8944 5280 8956
rect 5243 8436 5271 8944
rect 5234 8424 5280 8436
rect 5234 8390 5240 8424
rect 5274 8390 5280 8424
rect 5234 8378 5280 8390
rect 5243 8212 5271 8378
rect 5234 8200 5280 8212
rect 5234 8166 5240 8200
rect 5274 8166 5280 8200
rect 5234 8154 5280 8166
rect 5243 7646 5271 8154
rect 5234 7634 5280 7646
rect 5234 7600 5240 7634
rect 5274 7600 5280 7634
rect 5234 7588 5280 7600
rect 5243 7422 5271 7588
rect 5234 7410 5280 7422
rect 5234 7376 5240 7410
rect 5274 7376 5280 7410
rect 5234 7364 5280 7376
rect 5243 6856 5271 7364
rect 5234 6844 5280 6856
rect 5234 6810 5240 6844
rect 5274 6810 5280 6844
rect 5234 6798 5280 6810
rect 5243 6632 5271 6798
rect 5234 6620 5280 6632
rect 5234 6586 5240 6620
rect 5274 6586 5280 6620
rect 5234 6574 5280 6586
rect 5154 6054 5200 6066
rect 5154 6020 5160 6054
rect 5194 6020 5200 6054
rect 5154 6008 5200 6020
rect 5163 5842 5191 6008
rect 5154 5830 5200 5842
rect 5154 5796 5160 5830
rect 5194 5796 5200 5830
rect 5154 5784 5200 5796
rect 5074 5740 5120 5752
rect 5074 5706 5080 5740
rect 5114 5706 5120 5740
rect 5074 5694 5120 5706
rect 5083 5366 5111 5694
rect 5074 5354 5120 5366
rect 5074 5320 5080 5354
rect 5114 5320 5120 5354
rect 5074 5308 5120 5320
rect 5083 4962 5111 5308
rect 5163 5276 5191 5784
rect 5243 5332 5271 6574
rect 5323 5728 5351 12894
rect 5403 6122 5431 19214
rect 5483 6518 5511 25534
rect 5563 6912 5591 31854
rect 5643 7308 5671 38174
rect 5723 7702 5751 44494
rect 6051 44310 6097 44632
rect 6042 44258 6048 44310
rect 6100 44258 6106 44310
rect 6051 43894 6097 44258
rect 6475 44252 6523 44632
rect 6907 44252 6955 44632
rect 7281 44609 7287 44661
rect 7339 44609 7345 44661
rect 7677 44609 7683 44661
rect 7735 44609 7741 44661
rect 7299 44266 7327 44609
rect 7695 44266 7723 44609
rect 6467 44200 6473 44252
rect 6525 44200 6531 44252
rect 6899 44200 6905 44252
rect 6957 44200 6963 44252
rect 7281 44214 7287 44266
rect 7339 44214 7345 44266
rect 7677 44214 7683 44266
rect 7735 44214 7741 44266
rect 6475 43894 6523 44200
rect 6907 43894 6955 44200
rect 6042 43842 6048 43894
rect 6100 43842 6106 43894
rect 6467 43842 6473 43894
rect 6525 43842 6531 43894
rect 6899 43842 6905 43894
rect 6957 43842 6963 43894
rect 7299 43871 7327 44214
rect 7695 43871 7723 44214
rect 6051 43520 6097 43842
rect 6042 43468 6048 43520
rect 6100 43468 6106 43520
rect 6051 43104 6097 43468
rect 6475 43462 6523 43842
rect 6907 43462 6955 43842
rect 7281 43819 7287 43871
rect 7339 43819 7345 43871
rect 7677 43819 7683 43871
rect 7735 43819 7741 43871
rect 7299 43476 7327 43819
rect 7695 43476 7723 43819
rect 6467 43410 6473 43462
rect 6525 43410 6531 43462
rect 6899 43410 6905 43462
rect 6957 43410 6963 43462
rect 7281 43424 7287 43476
rect 7339 43424 7345 43476
rect 7677 43424 7683 43476
rect 7735 43424 7741 43476
rect 6475 43104 6523 43410
rect 6907 43104 6955 43410
rect 6042 43052 6048 43104
rect 6100 43052 6106 43104
rect 6467 43052 6473 43104
rect 6525 43052 6531 43104
rect 6899 43052 6905 43104
rect 6957 43052 6963 43104
rect 7299 43081 7327 43424
rect 7695 43081 7723 43424
rect 6051 42730 6097 43052
rect 6042 42678 6048 42730
rect 6100 42678 6106 42730
rect 6051 42314 6097 42678
rect 6475 42672 6523 43052
rect 6907 42672 6955 43052
rect 7281 43029 7287 43081
rect 7339 43029 7345 43081
rect 7677 43029 7683 43081
rect 7735 43029 7741 43081
rect 7299 42686 7327 43029
rect 7695 42686 7723 43029
rect 6467 42620 6473 42672
rect 6525 42620 6531 42672
rect 6899 42620 6905 42672
rect 6957 42620 6963 42672
rect 7281 42634 7287 42686
rect 7339 42634 7345 42686
rect 7677 42634 7683 42686
rect 7735 42634 7741 42686
rect 6475 42314 6523 42620
rect 6907 42314 6955 42620
rect 6042 42262 6048 42314
rect 6100 42262 6106 42314
rect 6467 42262 6473 42314
rect 6525 42262 6531 42314
rect 6899 42262 6905 42314
rect 6957 42262 6963 42314
rect 7299 42291 7327 42634
rect 7695 42291 7723 42634
rect 6051 41940 6097 42262
rect 6042 41888 6048 41940
rect 6100 41888 6106 41940
rect 6051 41524 6097 41888
rect 6475 41882 6523 42262
rect 6907 41882 6955 42262
rect 7281 42239 7287 42291
rect 7339 42239 7345 42291
rect 7677 42239 7683 42291
rect 7735 42239 7741 42291
rect 7299 41896 7327 42239
rect 7695 41896 7723 42239
rect 6467 41830 6473 41882
rect 6525 41830 6531 41882
rect 6899 41830 6905 41882
rect 6957 41830 6963 41882
rect 7281 41844 7287 41896
rect 7339 41844 7345 41896
rect 7677 41844 7683 41896
rect 7735 41844 7741 41896
rect 6475 41524 6523 41830
rect 6907 41524 6955 41830
rect 6042 41472 6048 41524
rect 6100 41472 6106 41524
rect 6467 41472 6473 41524
rect 6525 41472 6531 41524
rect 6899 41472 6905 41524
rect 6957 41472 6963 41524
rect 7299 41501 7327 41844
rect 7695 41501 7723 41844
rect 6051 41150 6097 41472
rect 6042 41098 6048 41150
rect 6100 41098 6106 41150
rect 6051 40734 6097 41098
rect 6475 41092 6523 41472
rect 6907 41092 6955 41472
rect 7281 41449 7287 41501
rect 7339 41449 7345 41501
rect 7677 41449 7683 41501
rect 7735 41449 7741 41501
rect 7299 41106 7327 41449
rect 7695 41106 7723 41449
rect 6467 41040 6473 41092
rect 6525 41040 6531 41092
rect 6899 41040 6905 41092
rect 6957 41040 6963 41092
rect 7281 41054 7287 41106
rect 7339 41054 7345 41106
rect 7677 41054 7683 41106
rect 7735 41054 7741 41106
rect 6475 40734 6523 41040
rect 6907 40734 6955 41040
rect 6042 40682 6048 40734
rect 6100 40682 6106 40734
rect 6467 40682 6473 40734
rect 6525 40682 6531 40734
rect 6899 40682 6905 40734
rect 6957 40682 6963 40734
rect 7299 40711 7327 41054
rect 7695 40711 7723 41054
rect 6051 40360 6097 40682
rect 6042 40308 6048 40360
rect 6100 40308 6106 40360
rect 6051 39944 6097 40308
rect 6475 40302 6523 40682
rect 6907 40302 6955 40682
rect 7281 40659 7287 40711
rect 7339 40659 7345 40711
rect 7677 40659 7683 40711
rect 7735 40659 7741 40711
rect 7299 40316 7327 40659
rect 7695 40316 7723 40659
rect 6467 40250 6473 40302
rect 6525 40250 6531 40302
rect 6899 40250 6905 40302
rect 6957 40250 6963 40302
rect 7281 40264 7287 40316
rect 7339 40264 7345 40316
rect 7677 40264 7683 40316
rect 7735 40264 7741 40316
rect 6475 39944 6523 40250
rect 6907 39944 6955 40250
rect 6042 39892 6048 39944
rect 6100 39892 6106 39944
rect 6467 39892 6473 39944
rect 6525 39892 6531 39944
rect 6899 39892 6905 39944
rect 6957 39892 6963 39944
rect 7299 39921 7327 40264
rect 7695 39921 7723 40264
rect 6051 39570 6097 39892
rect 6042 39518 6048 39570
rect 6100 39518 6106 39570
rect 6051 39154 6097 39518
rect 6475 39512 6523 39892
rect 6907 39512 6955 39892
rect 7281 39869 7287 39921
rect 7339 39869 7345 39921
rect 7677 39869 7683 39921
rect 7735 39869 7741 39921
rect 7299 39526 7327 39869
rect 7695 39526 7723 39869
rect 6467 39460 6473 39512
rect 6525 39460 6531 39512
rect 6899 39460 6905 39512
rect 6957 39460 6963 39512
rect 7281 39474 7287 39526
rect 7339 39474 7345 39526
rect 7677 39474 7683 39526
rect 7735 39474 7741 39526
rect 6475 39154 6523 39460
rect 6907 39154 6955 39460
rect 6042 39102 6048 39154
rect 6100 39102 6106 39154
rect 6467 39102 6473 39154
rect 6525 39102 6531 39154
rect 6899 39102 6905 39154
rect 6957 39102 6963 39154
rect 7299 39131 7327 39474
rect 7695 39131 7723 39474
rect 6051 38780 6097 39102
rect 6042 38728 6048 38780
rect 6100 38728 6106 38780
rect 6051 38364 6097 38728
rect 6475 38722 6523 39102
rect 6907 38722 6955 39102
rect 7281 39079 7287 39131
rect 7339 39079 7345 39131
rect 7677 39079 7683 39131
rect 7735 39079 7741 39131
rect 7299 38736 7327 39079
rect 7695 38736 7723 39079
rect 6467 38670 6473 38722
rect 6525 38670 6531 38722
rect 6899 38670 6905 38722
rect 6957 38670 6963 38722
rect 7281 38684 7287 38736
rect 7339 38684 7345 38736
rect 7677 38684 7683 38736
rect 7735 38684 7741 38736
rect 6475 38364 6523 38670
rect 6907 38364 6955 38670
rect 6042 38312 6048 38364
rect 6100 38312 6106 38364
rect 6467 38312 6473 38364
rect 6525 38312 6531 38364
rect 6899 38312 6905 38364
rect 6957 38312 6963 38364
rect 7299 38341 7327 38684
rect 7695 38341 7723 38684
rect 6051 37990 6097 38312
rect 6042 37938 6048 37990
rect 6100 37938 6106 37990
rect 6051 37574 6097 37938
rect 6475 37932 6523 38312
rect 6907 37932 6955 38312
rect 7281 38289 7287 38341
rect 7339 38289 7345 38341
rect 7677 38289 7683 38341
rect 7735 38289 7741 38341
rect 7299 37946 7327 38289
rect 7695 37946 7723 38289
rect 6467 37880 6473 37932
rect 6525 37880 6531 37932
rect 6899 37880 6905 37932
rect 6957 37880 6963 37932
rect 7281 37894 7287 37946
rect 7339 37894 7345 37946
rect 7677 37894 7683 37946
rect 7735 37894 7741 37946
rect 6475 37574 6523 37880
rect 6907 37574 6955 37880
rect 6042 37522 6048 37574
rect 6100 37522 6106 37574
rect 6467 37522 6473 37574
rect 6525 37522 6531 37574
rect 6899 37522 6905 37574
rect 6957 37522 6963 37574
rect 7299 37551 7327 37894
rect 7695 37551 7723 37894
rect 6051 37200 6097 37522
rect 6042 37148 6048 37200
rect 6100 37148 6106 37200
rect 6051 36784 6097 37148
rect 6475 37142 6523 37522
rect 6907 37142 6955 37522
rect 7281 37499 7287 37551
rect 7339 37499 7345 37551
rect 7677 37499 7683 37551
rect 7735 37499 7741 37551
rect 7299 37156 7327 37499
rect 7695 37156 7723 37499
rect 6467 37090 6473 37142
rect 6525 37090 6531 37142
rect 6899 37090 6905 37142
rect 6957 37090 6963 37142
rect 7281 37104 7287 37156
rect 7339 37104 7345 37156
rect 7677 37104 7683 37156
rect 7735 37104 7741 37156
rect 6475 36784 6523 37090
rect 6907 36784 6955 37090
rect 6042 36732 6048 36784
rect 6100 36732 6106 36784
rect 6467 36732 6473 36784
rect 6525 36732 6531 36784
rect 6899 36732 6905 36784
rect 6957 36732 6963 36784
rect 7299 36761 7327 37104
rect 7695 36761 7723 37104
rect 6051 36410 6097 36732
rect 6042 36358 6048 36410
rect 6100 36358 6106 36410
rect 6051 35994 6097 36358
rect 6475 36352 6523 36732
rect 6907 36352 6955 36732
rect 7281 36709 7287 36761
rect 7339 36709 7345 36761
rect 7677 36709 7683 36761
rect 7735 36709 7741 36761
rect 7299 36366 7327 36709
rect 7695 36366 7723 36709
rect 6467 36300 6473 36352
rect 6525 36300 6531 36352
rect 6899 36300 6905 36352
rect 6957 36300 6963 36352
rect 7281 36314 7287 36366
rect 7339 36314 7345 36366
rect 7677 36314 7683 36366
rect 7735 36314 7741 36366
rect 6475 35994 6523 36300
rect 6907 35994 6955 36300
rect 6042 35942 6048 35994
rect 6100 35942 6106 35994
rect 6467 35942 6473 35994
rect 6525 35942 6531 35994
rect 6899 35942 6905 35994
rect 6957 35942 6963 35994
rect 7299 35971 7327 36314
rect 7695 35971 7723 36314
rect 6051 35620 6097 35942
rect 6042 35568 6048 35620
rect 6100 35568 6106 35620
rect 6051 35204 6097 35568
rect 6475 35562 6523 35942
rect 6907 35562 6955 35942
rect 7281 35919 7287 35971
rect 7339 35919 7345 35971
rect 7677 35919 7683 35971
rect 7735 35919 7741 35971
rect 7299 35576 7327 35919
rect 7695 35576 7723 35919
rect 6467 35510 6473 35562
rect 6525 35510 6531 35562
rect 6899 35510 6905 35562
rect 6957 35510 6963 35562
rect 7281 35524 7287 35576
rect 7339 35524 7345 35576
rect 7677 35524 7683 35576
rect 7735 35524 7741 35576
rect 6475 35204 6523 35510
rect 6907 35204 6955 35510
rect 6042 35152 6048 35204
rect 6100 35152 6106 35204
rect 6467 35152 6473 35204
rect 6525 35152 6531 35204
rect 6899 35152 6905 35204
rect 6957 35152 6963 35204
rect 7299 35181 7327 35524
rect 7695 35181 7723 35524
rect 6051 34830 6097 35152
rect 6042 34778 6048 34830
rect 6100 34778 6106 34830
rect 6051 34414 6097 34778
rect 6475 34772 6523 35152
rect 6907 34772 6955 35152
rect 7281 35129 7287 35181
rect 7339 35129 7345 35181
rect 7677 35129 7683 35181
rect 7735 35129 7741 35181
rect 7299 34786 7327 35129
rect 7695 34786 7723 35129
rect 6467 34720 6473 34772
rect 6525 34720 6531 34772
rect 6899 34720 6905 34772
rect 6957 34720 6963 34772
rect 7281 34734 7287 34786
rect 7339 34734 7345 34786
rect 7677 34734 7683 34786
rect 7735 34734 7741 34786
rect 6475 34414 6523 34720
rect 6907 34414 6955 34720
rect 6042 34362 6048 34414
rect 6100 34362 6106 34414
rect 6467 34362 6473 34414
rect 6525 34362 6531 34414
rect 6899 34362 6905 34414
rect 6957 34362 6963 34414
rect 7299 34391 7327 34734
rect 7695 34391 7723 34734
rect 6051 34040 6097 34362
rect 6042 33988 6048 34040
rect 6100 33988 6106 34040
rect 6051 33624 6097 33988
rect 6475 33982 6523 34362
rect 6907 33982 6955 34362
rect 7281 34339 7287 34391
rect 7339 34339 7345 34391
rect 7677 34339 7683 34391
rect 7735 34339 7741 34391
rect 7299 33996 7327 34339
rect 7695 33996 7723 34339
rect 6467 33930 6473 33982
rect 6525 33930 6531 33982
rect 6899 33930 6905 33982
rect 6957 33930 6963 33982
rect 7281 33944 7287 33996
rect 7339 33944 7345 33996
rect 7677 33944 7683 33996
rect 7735 33944 7741 33996
rect 6475 33624 6523 33930
rect 6907 33624 6955 33930
rect 6042 33572 6048 33624
rect 6100 33572 6106 33624
rect 6467 33572 6473 33624
rect 6525 33572 6531 33624
rect 6899 33572 6905 33624
rect 6957 33572 6963 33624
rect 7299 33601 7327 33944
rect 7695 33601 7723 33944
rect 6051 33250 6097 33572
rect 6042 33198 6048 33250
rect 6100 33198 6106 33250
rect 6051 32834 6097 33198
rect 6475 33192 6523 33572
rect 6907 33192 6955 33572
rect 7281 33549 7287 33601
rect 7339 33549 7345 33601
rect 7677 33549 7683 33601
rect 7735 33549 7741 33601
rect 7299 33206 7327 33549
rect 7695 33206 7723 33549
rect 6467 33140 6473 33192
rect 6525 33140 6531 33192
rect 6899 33140 6905 33192
rect 6957 33140 6963 33192
rect 7281 33154 7287 33206
rect 7339 33154 7345 33206
rect 7677 33154 7683 33206
rect 7735 33154 7741 33206
rect 6475 32834 6523 33140
rect 6907 32834 6955 33140
rect 6042 32782 6048 32834
rect 6100 32782 6106 32834
rect 6467 32782 6473 32834
rect 6525 32782 6531 32834
rect 6899 32782 6905 32834
rect 6957 32782 6963 32834
rect 7299 32811 7327 33154
rect 7695 32811 7723 33154
rect 6051 32460 6097 32782
rect 6042 32408 6048 32460
rect 6100 32408 6106 32460
rect 6051 32044 6097 32408
rect 6475 32402 6523 32782
rect 6907 32402 6955 32782
rect 7281 32759 7287 32811
rect 7339 32759 7345 32811
rect 7677 32759 7683 32811
rect 7735 32759 7741 32811
rect 7299 32416 7327 32759
rect 7695 32416 7723 32759
rect 6467 32350 6473 32402
rect 6525 32350 6531 32402
rect 6899 32350 6905 32402
rect 6957 32350 6963 32402
rect 7281 32364 7287 32416
rect 7339 32364 7345 32416
rect 7677 32364 7683 32416
rect 7735 32364 7741 32416
rect 6475 32044 6523 32350
rect 6907 32044 6955 32350
rect 6042 31992 6048 32044
rect 6100 31992 6106 32044
rect 6467 31992 6473 32044
rect 6525 31992 6531 32044
rect 6899 31992 6905 32044
rect 6957 31992 6963 32044
rect 7299 32021 7327 32364
rect 7695 32021 7723 32364
rect 6051 31670 6097 31992
rect 6042 31618 6048 31670
rect 6100 31618 6106 31670
rect 6051 31254 6097 31618
rect 6475 31612 6523 31992
rect 6907 31612 6955 31992
rect 7281 31969 7287 32021
rect 7339 31969 7345 32021
rect 7677 31969 7683 32021
rect 7735 31969 7741 32021
rect 7299 31626 7327 31969
rect 7695 31626 7723 31969
rect 6467 31560 6473 31612
rect 6525 31560 6531 31612
rect 6899 31560 6905 31612
rect 6957 31560 6963 31612
rect 7281 31574 7287 31626
rect 7339 31574 7345 31626
rect 7677 31574 7683 31626
rect 7735 31574 7741 31626
rect 6475 31254 6523 31560
rect 6907 31254 6955 31560
rect 6042 31202 6048 31254
rect 6100 31202 6106 31254
rect 6467 31202 6473 31254
rect 6525 31202 6531 31254
rect 6899 31202 6905 31254
rect 6957 31202 6963 31254
rect 7299 31231 7327 31574
rect 7695 31231 7723 31574
rect 6051 30880 6097 31202
rect 6042 30828 6048 30880
rect 6100 30828 6106 30880
rect 6051 30464 6097 30828
rect 6475 30822 6523 31202
rect 6907 30822 6955 31202
rect 7281 31179 7287 31231
rect 7339 31179 7345 31231
rect 7677 31179 7683 31231
rect 7735 31179 7741 31231
rect 7299 30836 7327 31179
rect 7695 30836 7723 31179
rect 6467 30770 6473 30822
rect 6525 30770 6531 30822
rect 6899 30770 6905 30822
rect 6957 30770 6963 30822
rect 7281 30784 7287 30836
rect 7339 30784 7345 30836
rect 7677 30784 7683 30836
rect 7735 30784 7741 30836
rect 6475 30464 6523 30770
rect 6907 30464 6955 30770
rect 6042 30412 6048 30464
rect 6100 30412 6106 30464
rect 6467 30412 6473 30464
rect 6525 30412 6531 30464
rect 6899 30412 6905 30464
rect 6957 30412 6963 30464
rect 7299 30441 7327 30784
rect 7695 30441 7723 30784
rect 6051 30090 6097 30412
rect 6042 30038 6048 30090
rect 6100 30038 6106 30090
rect 6051 29674 6097 30038
rect 6475 30032 6523 30412
rect 6907 30032 6955 30412
rect 7281 30389 7287 30441
rect 7339 30389 7345 30441
rect 7677 30389 7683 30441
rect 7735 30389 7741 30441
rect 7299 30046 7327 30389
rect 7695 30046 7723 30389
rect 6467 29980 6473 30032
rect 6525 29980 6531 30032
rect 6899 29980 6905 30032
rect 6957 29980 6963 30032
rect 7281 29994 7287 30046
rect 7339 29994 7345 30046
rect 7677 29994 7683 30046
rect 7735 29994 7741 30046
rect 6475 29674 6523 29980
rect 6907 29674 6955 29980
rect 6042 29622 6048 29674
rect 6100 29622 6106 29674
rect 6467 29622 6473 29674
rect 6525 29622 6531 29674
rect 6899 29622 6905 29674
rect 6957 29622 6963 29674
rect 7299 29651 7327 29994
rect 7695 29651 7723 29994
rect 6051 29300 6097 29622
rect 6042 29248 6048 29300
rect 6100 29248 6106 29300
rect 6051 28884 6097 29248
rect 6475 29242 6523 29622
rect 6907 29242 6955 29622
rect 7281 29599 7287 29651
rect 7339 29599 7345 29651
rect 7677 29599 7683 29651
rect 7735 29599 7741 29651
rect 7299 29256 7327 29599
rect 7695 29256 7723 29599
rect 6467 29190 6473 29242
rect 6525 29190 6531 29242
rect 6899 29190 6905 29242
rect 6957 29190 6963 29242
rect 7281 29204 7287 29256
rect 7339 29204 7345 29256
rect 7677 29204 7683 29256
rect 7735 29204 7741 29256
rect 6475 28884 6523 29190
rect 6907 28884 6955 29190
rect 6042 28832 6048 28884
rect 6100 28832 6106 28884
rect 6467 28832 6473 28884
rect 6525 28832 6531 28884
rect 6899 28832 6905 28884
rect 6957 28832 6963 28884
rect 7299 28861 7327 29204
rect 7695 28861 7723 29204
rect 6051 28510 6097 28832
rect 6042 28458 6048 28510
rect 6100 28458 6106 28510
rect 6051 28094 6097 28458
rect 6475 28452 6523 28832
rect 6907 28452 6955 28832
rect 7281 28809 7287 28861
rect 7339 28809 7345 28861
rect 7677 28809 7683 28861
rect 7735 28809 7741 28861
rect 7299 28466 7327 28809
rect 7695 28466 7723 28809
rect 6467 28400 6473 28452
rect 6525 28400 6531 28452
rect 6899 28400 6905 28452
rect 6957 28400 6963 28452
rect 7281 28414 7287 28466
rect 7339 28414 7345 28466
rect 7677 28414 7683 28466
rect 7735 28414 7741 28466
rect 6475 28094 6523 28400
rect 6907 28094 6955 28400
rect 6042 28042 6048 28094
rect 6100 28042 6106 28094
rect 6467 28042 6473 28094
rect 6525 28042 6531 28094
rect 6899 28042 6905 28094
rect 6957 28042 6963 28094
rect 7299 28071 7327 28414
rect 7695 28071 7723 28414
rect 6051 27720 6097 28042
rect 6042 27668 6048 27720
rect 6100 27668 6106 27720
rect 6051 27304 6097 27668
rect 6475 27662 6523 28042
rect 6907 27662 6955 28042
rect 7281 28019 7287 28071
rect 7339 28019 7345 28071
rect 7677 28019 7683 28071
rect 7735 28019 7741 28071
rect 7299 27676 7327 28019
rect 7695 27676 7723 28019
rect 6467 27610 6473 27662
rect 6525 27610 6531 27662
rect 6899 27610 6905 27662
rect 6957 27610 6963 27662
rect 7281 27624 7287 27676
rect 7339 27624 7345 27676
rect 7677 27624 7683 27676
rect 7735 27624 7741 27676
rect 6475 27304 6523 27610
rect 6907 27304 6955 27610
rect 6042 27252 6048 27304
rect 6100 27252 6106 27304
rect 6467 27252 6473 27304
rect 6525 27252 6531 27304
rect 6899 27252 6905 27304
rect 6957 27252 6963 27304
rect 7299 27281 7327 27624
rect 7695 27281 7723 27624
rect 6051 26930 6097 27252
rect 6042 26878 6048 26930
rect 6100 26878 6106 26930
rect 6051 26514 6097 26878
rect 6475 26872 6523 27252
rect 6907 26872 6955 27252
rect 7281 27229 7287 27281
rect 7339 27229 7345 27281
rect 7677 27229 7683 27281
rect 7735 27229 7741 27281
rect 7299 26886 7327 27229
rect 7695 26886 7723 27229
rect 6467 26820 6473 26872
rect 6525 26820 6531 26872
rect 6899 26820 6905 26872
rect 6957 26820 6963 26872
rect 7281 26834 7287 26886
rect 7339 26834 7345 26886
rect 7677 26834 7683 26886
rect 7735 26834 7741 26886
rect 6475 26514 6523 26820
rect 6907 26514 6955 26820
rect 6042 26462 6048 26514
rect 6100 26462 6106 26514
rect 6467 26462 6473 26514
rect 6525 26462 6531 26514
rect 6899 26462 6905 26514
rect 6957 26462 6963 26514
rect 7299 26491 7327 26834
rect 7695 26491 7723 26834
rect 6051 26140 6097 26462
rect 6042 26088 6048 26140
rect 6100 26088 6106 26140
rect 6051 25724 6097 26088
rect 6475 26082 6523 26462
rect 6907 26082 6955 26462
rect 7281 26439 7287 26491
rect 7339 26439 7345 26491
rect 7677 26439 7683 26491
rect 7735 26439 7741 26491
rect 7299 26096 7327 26439
rect 7695 26096 7723 26439
rect 6467 26030 6473 26082
rect 6525 26030 6531 26082
rect 6899 26030 6905 26082
rect 6957 26030 6963 26082
rect 7281 26044 7287 26096
rect 7339 26044 7345 26096
rect 7677 26044 7683 26096
rect 7735 26044 7741 26096
rect 6475 25724 6523 26030
rect 6907 25724 6955 26030
rect 6042 25672 6048 25724
rect 6100 25672 6106 25724
rect 6467 25672 6473 25724
rect 6525 25672 6531 25724
rect 6899 25672 6905 25724
rect 6957 25672 6963 25724
rect 7299 25701 7327 26044
rect 7695 25701 7723 26044
rect 6051 25350 6097 25672
rect 6042 25298 6048 25350
rect 6100 25298 6106 25350
rect 6051 24934 6097 25298
rect 6475 25292 6523 25672
rect 6907 25292 6955 25672
rect 7281 25649 7287 25701
rect 7339 25649 7345 25701
rect 7677 25649 7683 25701
rect 7735 25649 7741 25701
rect 7299 25306 7327 25649
rect 7695 25306 7723 25649
rect 6467 25240 6473 25292
rect 6525 25240 6531 25292
rect 6899 25240 6905 25292
rect 6957 25240 6963 25292
rect 7281 25254 7287 25306
rect 7339 25254 7345 25306
rect 7677 25254 7683 25306
rect 7735 25254 7741 25306
rect 6475 24934 6523 25240
rect 6907 24934 6955 25240
rect 6042 24882 6048 24934
rect 6100 24882 6106 24934
rect 6467 24882 6473 24934
rect 6525 24882 6531 24934
rect 6899 24882 6905 24934
rect 6957 24882 6963 24934
rect 7299 24911 7327 25254
rect 7695 24911 7723 25254
rect 6051 24560 6097 24882
rect 6042 24508 6048 24560
rect 6100 24508 6106 24560
rect 6051 24144 6097 24508
rect 6475 24502 6523 24882
rect 6907 24502 6955 24882
rect 7281 24859 7287 24911
rect 7339 24859 7345 24911
rect 7677 24859 7683 24911
rect 7735 24859 7741 24911
rect 7299 24516 7327 24859
rect 7695 24516 7723 24859
rect 6467 24450 6473 24502
rect 6525 24450 6531 24502
rect 6899 24450 6905 24502
rect 6957 24450 6963 24502
rect 7281 24464 7287 24516
rect 7339 24464 7345 24516
rect 7677 24464 7683 24516
rect 7735 24464 7741 24516
rect 6475 24144 6523 24450
rect 6907 24144 6955 24450
rect 6042 24092 6048 24144
rect 6100 24092 6106 24144
rect 6467 24092 6473 24144
rect 6525 24092 6531 24144
rect 6899 24092 6905 24144
rect 6957 24092 6963 24144
rect 7299 24121 7327 24464
rect 7695 24121 7723 24464
rect 6051 23770 6097 24092
rect 6042 23718 6048 23770
rect 6100 23718 6106 23770
rect 6051 23354 6097 23718
rect 6475 23712 6523 24092
rect 6907 23712 6955 24092
rect 7281 24069 7287 24121
rect 7339 24069 7345 24121
rect 7677 24069 7683 24121
rect 7735 24069 7741 24121
rect 7299 23726 7327 24069
rect 7695 23726 7723 24069
rect 6467 23660 6473 23712
rect 6525 23660 6531 23712
rect 6899 23660 6905 23712
rect 6957 23660 6963 23712
rect 7281 23674 7287 23726
rect 7339 23674 7345 23726
rect 7677 23674 7683 23726
rect 7735 23674 7741 23726
rect 6475 23354 6523 23660
rect 6907 23354 6955 23660
rect 6042 23302 6048 23354
rect 6100 23302 6106 23354
rect 6467 23302 6473 23354
rect 6525 23302 6531 23354
rect 6899 23302 6905 23354
rect 6957 23302 6963 23354
rect 7299 23331 7327 23674
rect 7695 23331 7723 23674
rect 6051 22980 6097 23302
rect 6042 22928 6048 22980
rect 6100 22928 6106 22980
rect 6051 22564 6097 22928
rect 6475 22922 6523 23302
rect 6907 22922 6955 23302
rect 7281 23279 7287 23331
rect 7339 23279 7345 23331
rect 7677 23279 7683 23331
rect 7735 23279 7741 23331
rect 7299 22936 7327 23279
rect 7695 22936 7723 23279
rect 6467 22870 6473 22922
rect 6525 22870 6531 22922
rect 6899 22870 6905 22922
rect 6957 22870 6963 22922
rect 7281 22884 7287 22936
rect 7339 22884 7345 22936
rect 7677 22884 7683 22936
rect 7735 22884 7741 22936
rect 6475 22564 6523 22870
rect 6907 22564 6955 22870
rect 6042 22512 6048 22564
rect 6100 22512 6106 22564
rect 6467 22512 6473 22564
rect 6525 22512 6531 22564
rect 6899 22512 6905 22564
rect 6957 22512 6963 22564
rect 7299 22541 7327 22884
rect 7695 22541 7723 22884
rect 6051 22190 6097 22512
rect 6042 22138 6048 22190
rect 6100 22138 6106 22190
rect 6051 21774 6097 22138
rect 6475 22132 6523 22512
rect 6907 22132 6955 22512
rect 7281 22489 7287 22541
rect 7339 22489 7345 22541
rect 7677 22489 7683 22541
rect 7735 22489 7741 22541
rect 7299 22146 7327 22489
rect 7695 22146 7723 22489
rect 6467 22080 6473 22132
rect 6525 22080 6531 22132
rect 6899 22080 6905 22132
rect 6957 22080 6963 22132
rect 7281 22094 7287 22146
rect 7339 22094 7345 22146
rect 7677 22094 7683 22146
rect 7735 22094 7741 22146
rect 6475 21774 6523 22080
rect 6907 21774 6955 22080
rect 6042 21722 6048 21774
rect 6100 21722 6106 21774
rect 6467 21722 6473 21774
rect 6525 21722 6531 21774
rect 6899 21722 6905 21774
rect 6957 21722 6963 21774
rect 7299 21751 7327 22094
rect 7695 21751 7723 22094
rect 6051 21400 6097 21722
rect 6042 21348 6048 21400
rect 6100 21348 6106 21400
rect 6051 20984 6097 21348
rect 6475 21342 6523 21722
rect 6907 21342 6955 21722
rect 7281 21699 7287 21751
rect 7339 21699 7345 21751
rect 7677 21699 7683 21751
rect 7735 21699 7741 21751
rect 7299 21356 7327 21699
rect 7695 21356 7723 21699
rect 6467 21290 6473 21342
rect 6525 21290 6531 21342
rect 6899 21290 6905 21342
rect 6957 21290 6963 21342
rect 7281 21304 7287 21356
rect 7339 21304 7345 21356
rect 7677 21304 7683 21356
rect 7735 21304 7741 21356
rect 6475 20984 6523 21290
rect 6907 20984 6955 21290
rect 6042 20932 6048 20984
rect 6100 20932 6106 20984
rect 6467 20932 6473 20984
rect 6525 20932 6531 20984
rect 6899 20932 6905 20984
rect 6957 20932 6963 20984
rect 7299 20961 7327 21304
rect 7695 20961 7723 21304
rect 6051 20610 6097 20932
rect 6042 20558 6048 20610
rect 6100 20558 6106 20610
rect 6051 20194 6097 20558
rect 6475 20552 6523 20932
rect 6907 20552 6955 20932
rect 7281 20909 7287 20961
rect 7339 20909 7345 20961
rect 7677 20909 7683 20961
rect 7735 20909 7741 20961
rect 7299 20566 7327 20909
rect 7695 20566 7723 20909
rect 6467 20500 6473 20552
rect 6525 20500 6531 20552
rect 6899 20500 6905 20552
rect 6957 20500 6963 20552
rect 7281 20514 7287 20566
rect 7339 20514 7345 20566
rect 7677 20514 7683 20566
rect 7735 20514 7741 20566
rect 6475 20194 6523 20500
rect 6907 20194 6955 20500
rect 6042 20142 6048 20194
rect 6100 20142 6106 20194
rect 6467 20142 6473 20194
rect 6525 20142 6531 20194
rect 6899 20142 6905 20194
rect 6957 20142 6963 20194
rect 7299 20171 7327 20514
rect 7695 20171 7723 20514
rect 6051 19820 6097 20142
rect 6042 19768 6048 19820
rect 6100 19768 6106 19820
rect 6051 19404 6097 19768
rect 6475 19762 6523 20142
rect 6907 19762 6955 20142
rect 7281 20119 7287 20171
rect 7339 20119 7345 20171
rect 7677 20119 7683 20171
rect 7735 20119 7741 20171
rect 7299 19776 7327 20119
rect 7695 19776 7723 20119
rect 6467 19710 6473 19762
rect 6525 19710 6531 19762
rect 6899 19710 6905 19762
rect 6957 19710 6963 19762
rect 7281 19724 7287 19776
rect 7339 19724 7345 19776
rect 7677 19724 7683 19776
rect 7735 19724 7741 19776
rect 6475 19404 6523 19710
rect 6907 19404 6955 19710
rect 6042 19352 6048 19404
rect 6100 19352 6106 19404
rect 6467 19352 6473 19404
rect 6525 19352 6531 19404
rect 6899 19352 6905 19404
rect 6957 19352 6963 19404
rect 7299 19381 7327 19724
rect 7695 19381 7723 19724
rect 6051 19030 6097 19352
rect 6042 18978 6048 19030
rect 6100 18978 6106 19030
rect 6051 18614 6097 18978
rect 6475 18972 6523 19352
rect 6907 18972 6955 19352
rect 7281 19329 7287 19381
rect 7339 19329 7345 19381
rect 7677 19329 7683 19381
rect 7735 19329 7741 19381
rect 7299 18986 7327 19329
rect 7695 18986 7723 19329
rect 6467 18920 6473 18972
rect 6525 18920 6531 18972
rect 6899 18920 6905 18972
rect 6957 18920 6963 18972
rect 7281 18934 7287 18986
rect 7339 18934 7345 18986
rect 7677 18934 7683 18986
rect 7735 18934 7741 18986
rect 6475 18614 6523 18920
rect 6907 18614 6955 18920
rect 6042 18562 6048 18614
rect 6100 18562 6106 18614
rect 6467 18562 6473 18614
rect 6525 18562 6531 18614
rect 6899 18562 6905 18614
rect 6957 18562 6963 18614
rect 7299 18591 7327 18934
rect 7695 18591 7723 18934
rect 6051 18240 6097 18562
rect 6042 18188 6048 18240
rect 6100 18188 6106 18240
rect 6051 17824 6097 18188
rect 6475 18182 6523 18562
rect 6907 18182 6955 18562
rect 7281 18539 7287 18591
rect 7339 18539 7345 18591
rect 7677 18539 7683 18591
rect 7735 18539 7741 18591
rect 7299 18196 7327 18539
rect 7695 18196 7723 18539
rect 6467 18130 6473 18182
rect 6525 18130 6531 18182
rect 6899 18130 6905 18182
rect 6957 18130 6963 18182
rect 7281 18144 7287 18196
rect 7339 18144 7345 18196
rect 7677 18144 7683 18196
rect 7735 18144 7741 18196
rect 6475 17824 6523 18130
rect 6907 17824 6955 18130
rect 6042 17772 6048 17824
rect 6100 17772 6106 17824
rect 6467 17772 6473 17824
rect 6525 17772 6531 17824
rect 6899 17772 6905 17824
rect 6957 17772 6963 17824
rect 7299 17801 7327 18144
rect 7695 17801 7723 18144
rect 6051 17450 6097 17772
rect 6042 17398 6048 17450
rect 6100 17398 6106 17450
rect 6051 17034 6097 17398
rect 6475 17392 6523 17772
rect 6907 17392 6955 17772
rect 7281 17749 7287 17801
rect 7339 17749 7345 17801
rect 7677 17749 7683 17801
rect 7735 17749 7741 17801
rect 7299 17406 7327 17749
rect 7695 17406 7723 17749
rect 6467 17340 6473 17392
rect 6525 17340 6531 17392
rect 6899 17340 6905 17392
rect 6957 17340 6963 17392
rect 7281 17354 7287 17406
rect 7339 17354 7345 17406
rect 7677 17354 7683 17406
rect 7735 17354 7741 17406
rect 6475 17034 6523 17340
rect 6907 17034 6955 17340
rect 6042 16982 6048 17034
rect 6100 16982 6106 17034
rect 6467 16982 6473 17034
rect 6525 16982 6531 17034
rect 6899 16982 6905 17034
rect 6957 16982 6963 17034
rect 7299 17011 7327 17354
rect 7695 17011 7723 17354
rect 6051 16660 6097 16982
rect 6042 16608 6048 16660
rect 6100 16608 6106 16660
rect 6051 16244 6097 16608
rect 6475 16602 6523 16982
rect 6907 16602 6955 16982
rect 7281 16959 7287 17011
rect 7339 16959 7345 17011
rect 7677 16959 7683 17011
rect 7735 16959 7741 17011
rect 7299 16616 7327 16959
rect 7695 16616 7723 16959
rect 6467 16550 6473 16602
rect 6525 16550 6531 16602
rect 6899 16550 6905 16602
rect 6957 16550 6963 16602
rect 7281 16564 7287 16616
rect 7339 16564 7345 16616
rect 7677 16564 7683 16616
rect 7735 16564 7741 16616
rect 6475 16244 6523 16550
rect 6907 16244 6955 16550
rect 6042 16192 6048 16244
rect 6100 16192 6106 16244
rect 6467 16192 6473 16244
rect 6525 16192 6531 16244
rect 6899 16192 6905 16244
rect 6957 16192 6963 16244
rect 7299 16221 7327 16564
rect 7695 16221 7723 16564
rect 6051 15870 6097 16192
rect 6042 15818 6048 15870
rect 6100 15818 6106 15870
rect 6051 15454 6097 15818
rect 6475 15812 6523 16192
rect 6907 15812 6955 16192
rect 7281 16169 7287 16221
rect 7339 16169 7345 16221
rect 7677 16169 7683 16221
rect 7735 16169 7741 16221
rect 7299 15826 7327 16169
rect 7695 15826 7723 16169
rect 6467 15760 6473 15812
rect 6525 15760 6531 15812
rect 6899 15760 6905 15812
rect 6957 15760 6963 15812
rect 7281 15774 7287 15826
rect 7339 15774 7345 15826
rect 7677 15774 7683 15826
rect 7735 15774 7741 15826
rect 6475 15454 6523 15760
rect 6907 15454 6955 15760
rect 6042 15402 6048 15454
rect 6100 15402 6106 15454
rect 6467 15402 6473 15454
rect 6525 15402 6531 15454
rect 6899 15402 6905 15454
rect 6957 15402 6963 15454
rect 7299 15431 7327 15774
rect 7695 15431 7723 15774
rect 6051 15080 6097 15402
rect 6042 15028 6048 15080
rect 6100 15028 6106 15080
rect 6051 14664 6097 15028
rect 6475 15022 6523 15402
rect 6907 15022 6955 15402
rect 7281 15379 7287 15431
rect 7339 15379 7345 15431
rect 7677 15379 7683 15431
rect 7735 15379 7741 15431
rect 7299 15036 7327 15379
rect 7695 15036 7723 15379
rect 6467 14970 6473 15022
rect 6525 14970 6531 15022
rect 6899 14970 6905 15022
rect 6957 14970 6963 15022
rect 7281 14984 7287 15036
rect 7339 14984 7345 15036
rect 7677 14984 7683 15036
rect 7735 14984 7741 15036
rect 6475 14664 6523 14970
rect 6907 14664 6955 14970
rect 6042 14612 6048 14664
rect 6100 14612 6106 14664
rect 6467 14612 6473 14664
rect 6525 14612 6531 14664
rect 6899 14612 6905 14664
rect 6957 14612 6963 14664
rect 7299 14641 7327 14984
rect 7695 14641 7723 14984
rect 6051 14290 6097 14612
rect 6042 14238 6048 14290
rect 6100 14238 6106 14290
rect 6051 13874 6097 14238
rect 6475 14232 6523 14612
rect 6907 14232 6955 14612
rect 7281 14589 7287 14641
rect 7339 14589 7345 14641
rect 7677 14589 7683 14641
rect 7735 14589 7741 14641
rect 7299 14246 7327 14589
rect 7695 14246 7723 14589
rect 6467 14180 6473 14232
rect 6525 14180 6531 14232
rect 6899 14180 6905 14232
rect 6957 14180 6963 14232
rect 7281 14194 7287 14246
rect 7339 14194 7345 14246
rect 7677 14194 7683 14246
rect 7735 14194 7741 14246
rect 6475 13874 6523 14180
rect 6907 13874 6955 14180
rect 6042 13822 6048 13874
rect 6100 13822 6106 13874
rect 6467 13822 6473 13874
rect 6525 13822 6531 13874
rect 6899 13822 6905 13874
rect 6957 13822 6963 13874
rect 7299 13851 7327 14194
rect 7695 13851 7723 14194
rect 6051 13500 6097 13822
rect 6042 13448 6048 13500
rect 6100 13448 6106 13500
rect 6051 13084 6097 13448
rect 6475 13442 6523 13822
rect 6907 13442 6955 13822
rect 7281 13799 7287 13851
rect 7339 13799 7345 13851
rect 7677 13799 7683 13851
rect 7735 13799 7741 13851
rect 7299 13456 7327 13799
rect 7695 13456 7723 13799
rect 6467 13390 6473 13442
rect 6525 13390 6531 13442
rect 6899 13390 6905 13442
rect 6957 13390 6963 13442
rect 7281 13404 7287 13456
rect 7339 13404 7345 13456
rect 7677 13404 7683 13456
rect 7735 13404 7741 13456
rect 6475 13084 6523 13390
rect 6907 13084 6955 13390
rect 6042 13032 6048 13084
rect 6100 13032 6106 13084
rect 6467 13032 6473 13084
rect 6525 13032 6531 13084
rect 6899 13032 6905 13084
rect 6957 13032 6963 13084
rect 7299 13061 7327 13404
rect 7695 13061 7723 13404
rect 6051 12710 6097 13032
rect 6042 12658 6048 12710
rect 6100 12658 6106 12710
rect 6051 12294 6097 12658
rect 6475 12652 6523 13032
rect 6907 12652 6955 13032
rect 7281 13009 7287 13061
rect 7339 13009 7345 13061
rect 7677 13009 7683 13061
rect 7735 13009 7741 13061
rect 7299 12666 7327 13009
rect 7695 12666 7723 13009
rect 6467 12600 6473 12652
rect 6525 12600 6531 12652
rect 6899 12600 6905 12652
rect 6957 12600 6963 12652
rect 7281 12614 7287 12666
rect 7339 12614 7345 12666
rect 7677 12614 7683 12666
rect 7735 12614 7741 12666
rect 6475 12294 6523 12600
rect 6907 12294 6955 12600
rect 6042 12242 6048 12294
rect 6100 12242 6106 12294
rect 6467 12242 6473 12294
rect 6525 12242 6531 12294
rect 6899 12242 6905 12294
rect 6957 12242 6963 12294
rect 7299 12271 7327 12614
rect 7695 12271 7723 12614
rect 6051 11920 6097 12242
rect 6042 11868 6048 11920
rect 6100 11868 6106 11920
rect 6051 11504 6097 11868
rect 6475 11862 6523 12242
rect 6907 11862 6955 12242
rect 7281 12219 7287 12271
rect 7339 12219 7345 12271
rect 7677 12219 7683 12271
rect 7735 12219 7741 12271
rect 7299 11876 7327 12219
rect 7695 11876 7723 12219
rect 6467 11810 6473 11862
rect 6525 11810 6531 11862
rect 6899 11810 6905 11862
rect 6957 11810 6963 11862
rect 7281 11824 7287 11876
rect 7339 11824 7345 11876
rect 7677 11824 7683 11876
rect 7735 11824 7741 11876
rect 6475 11504 6523 11810
rect 6907 11504 6955 11810
rect 6042 11452 6048 11504
rect 6100 11452 6106 11504
rect 6467 11452 6473 11504
rect 6525 11452 6531 11504
rect 6899 11452 6905 11504
rect 6957 11452 6963 11504
rect 7299 11481 7327 11824
rect 7695 11481 7723 11824
rect 6051 11130 6097 11452
rect 6042 11078 6048 11130
rect 6100 11078 6106 11130
rect 6051 10714 6097 11078
rect 6475 11072 6523 11452
rect 6907 11072 6955 11452
rect 7281 11429 7287 11481
rect 7339 11429 7345 11481
rect 7677 11429 7683 11481
rect 7735 11429 7741 11481
rect 7299 11086 7327 11429
rect 7695 11086 7723 11429
rect 6467 11020 6473 11072
rect 6525 11020 6531 11072
rect 6899 11020 6905 11072
rect 6957 11020 6963 11072
rect 7281 11034 7287 11086
rect 7339 11034 7345 11086
rect 7677 11034 7683 11086
rect 7735 11034 7741 11086
rect 6475 10714 6523 11020
rect 6907 10714 6955 11020
rect 6042 10662 6048 10714
rect 6100 10662 6106 10714
rect 6467 10662 6473 10714
rect 6525 10662 6531 10714
rect 6899 10662 6905 10714
rect 6957 10662 6963 10714
rect 7299 10691 7327 11034
rect 7695 10691 7723 11034
rect 6051 10340 6097 10662
rect 6042 10288 6048 10340
rect 6100 10288 6106 10340
rect 6051 9924 6097 10288
rect 6475 10282 6523 10662
rect 6907 10282 6955 10662
rect 7281 10639 7287 10691
rect 7339 10639 7345 10691
rect 7677 10639 7683 10691
rect 7735 10639 7741 10691
rect 7299 10296 7327 10639
rect 7695 10296 7723 10639
rect 6467 10230 6473 10282
rect 6525 10230 6531 10282
rect 6899 10230 6905 10282
rect 6957 10230 6963 10282
rect 7281 10244 7287 10296
rect 7339 10244 7345 10296
rect 7677 10244 7683 10296
rect 7735 10244 7741 10296
rect 6475 9924 6523 10230
rect 6907 9924 6955 10230
rect 6042 9872 6048 9924
rect 6100 9872 6106 9924
rect 6467 9872 6473 9924
rect 6525 9872 6531 9924
rect 6899 9872 6905 9924
rect 6957 9872 6963 9924
rect 7299 9901 7327 10244
rect 7695 9901 7723 10244
rect 6051 9550 6097 9872
rect 6042 9498 6048 9550
rect 6100 9498 6106 9550
rect 6051 9134 6097 9498
rect 6475 9492 6523 9872
rect 6907 9492 6955 9872
rect 7281 9849 7287 9901
rect 7339 9849 7345 9901
rect 7677 9849 7683 9901
rect 7735 9849 7741 9901
rect 7299 9506 7327 9849
rect 7695 9506 7723 9849
rect 6467 9440 6473 9492
rect 6525 9440 6531 9492
rect 6899 9440 6905 9492
rect 6957 9440 6963 9492
rect 7281 9454 7287 9506
rect 7339 9454 7345 9506
rect 7677 9454 7683 9506
rect 7735 9454 7741 9506
rect 6475 9134 6523 9440
rect 6907 9134 6955 9440
rect 6042 9082 6048 9134
rect 6100 9082 6106 9134
rect 6467 9082 6473 9134
rect 6525 9082 6531 9134
rect 6899 9082 6905 9134
rect 6957 9082 6963 9134
rect 7299 9111 7327 9454
rect 7695 9111 7723 9454
rect 6051 8760 6097 9082
rect 6042 8708 6048 8760
rect 6100 8708 6106 8760
rect 6051 8344 6097 8708
rect 6475 8702 6523 9082
rect 6907 8702 6955 9082
rect 7281 9059 7287 9111
rect 7339 9059 7345 9111
rect 7677 9059 7683 9111
rect 7735 9059 7741 9111
rect 7299 8716 7327 9059
rect 7695 8716 7723 9059
rect 6467 8650 6473 8702
rect 6525 8650 6531 8702
rect 6899 8650 6905 8702
rect 6957 8650 6963 8702
rect 7281 8664 7287 8716
rect 7339 8664 7345 8716
rect 7677 8664 7683 8716
rect 7735 8664 7741 8716
rect 6475 8344 6523 8650
rect 6907 8344 6955 8650
rect 6042 8292 6048 8344
rect 6100 8292 6106 8344
rect 6467 8292 6473 8344
rect 6525 8292 6531 8344
rect 6899 8292 6905 8344
rect 6957 8292 6963 8344
rect 7299 8321 7327 8664
rect 7695 8321 7723 8664
rect 6051 7970 6097 8292
rect 6042 7918 6048 7970
rect 6100 7918 6106 7970
rect 5714 7537 5760 7702
rect 6051 7554 6097 7918
rect 6475 7912 6523 8292
rect 6907 7912 6955 8292
rect 7281 8269 7287 8321
rect 7339 8269 7345 8321
rect 7677 8269 7683 8321
rect 7735 8269 7741 8321
rect 7299 7926 7327 8269
rect 7695 7926 7723 8269
rect 6467 7860 6473 7912
rect 6525 7860 6531 7912
rect 6899 7860 6905 7912
rect 6957 7860 6963 7912
rect 7281 7874 7287 7926
rect 7339 7874 7345 7926
rect 7677 7874 7683 7926
rect 7735 7874 7741 7926
rect 6475 7554 6523 7860
rect 6907 7554 6955 7860
rect 5711 7531 5763 7537
rect 6042 7502 6048 7554
rect 6100 7502 6106 7554
rect 6467 7502 6473 7554
rect 6525 7502 6531 7554
rect 6899 7502 6905 7554
rect 6957 7502 6963 7554
rect 7299 7531 7327 7874
rect 7695 7531 7723 7874
rect 5711 7473 5763 7479
rect 5634 7142 5680 7308
rect 5631 7136 5683 7142
rect 5631 7078 5683 7084
rect 5554 6747 5600 6912
rect 5551 6741 5603 6747
rect 5551 6683 5603 6689
rect 5474 6352 5520 6518
rect 5471 6346 5523 6352
rect 5471 6288 5523 6294
rect 5394 5957 5440 6122
rect 5391 5951 5443 5957
rect 5391 5893 5443 5899
rect 5314 5562 5360 5728
rect 5311 5556 5363 5562
rect 5311 5498 5363 5504
rect 5154 5264 5200 5276
rect 5154 5230 5160 5264
rect 5194 5230 5200 5264
rect 5154 5218 5200 5230
rect 5163 5052 5191 5218
rect 5234 5167 5280 5332
rect 5231 5161 5283 5167
rect 5231 5103 5283 5109
rect 5154 5040 5200 5052
rect 5154 5006 5160 5040
rect 5194 5006 5200 5040
rect 5154 4994 5200 5006
rect 5074 4950 5120 4962
rect 5074 4916 5080 4950
rect 5114 4916 5120 4950
rect 5163 4938 5191 4994
rect 5074 4904 5120 4916
rect 4994 4564 5040 4576
rect 4994 4530 5000 4564
rect 5034 4530 5040 4564
rect 4994 4518 5040 4530
rect 5003 4172 5031 4518
rect 4994 4160 5040 4172
rect 4994 4126 5000 4160
rect 5034 4126 5040 4160
rect 4994 4114 5040 4126
rect 5003 3786 5031 4114
rect 4994 3774 5040 3786
rect 4994 3740 5000 3774
rect 5034 3740 5040 3774
rect 5083 3752 5111 4904
rect 5154 4772 5200 4938
rect 5151 4766 5203 4772
rect 5151 4708 5203 4714
rect 5163 4486 5191 4708
rect 5154 4474 5200 4486
rect 5154 4440 5160 4474
rect 5194 4440 5200 4474
rect 5154 4428 5200 4440
rect 5163 4262 5191 4428
rect 5154 4250 5200 4262
rect 5154 4216 5160 4250
rect 5194 4216 5200 4250
rect 5154 4204 5200 4216
rect 4994 3728 5040 3740
rect 5003 3382 5031 3728
rect 5074 3587 5120 3752
rect 5163 3696 5191 4204
rect 5154 3684 5200 3696
rect 5154 3650 5160 3684
rect 5194 3650 5200 3684
rect 5154 3638 5200 3650
rect 5071 3581 5123 3587
rect 5071 3523 5123 3529
rect 4994 3370 5040 3382
rect 4994 3336 5000 3370
rect 5034 3336 5040 3370
rect 4994 3192 5040 3336
rect 4991 3186 5043 3192
rect 4991 3128 5043 3134
rect 4914 2984 4960 2996
rect 4914 2950 4920 2984
rect 4954 2950 4960 2984
rect 4914 2797 4960 2950
rect 4911 2791 4963 2797
rect 4911 2733 4963 2739
rect 4923 2592 4951 2733
rect 4914 2580 4960 2592
rect 4834 2402 4880 2568
rect 4914 2546 4920 2580
rect 4954 2546 4960 2580
rect 4914 2534 4960 2546
rect 4831 2396 4883 2402
rect 4831 2338 4883 2344
rect 4754 1516 4800 1528
rect 4754 1482 4760 1516
rect 4794 1482 4800 1516
rect 4754 1470 4800 1482
rect 4763 1382 4791 1470
rect 4843 1416 4871 2338
rect 4923 2206 4951 2534
rect 4914 2194 4960 2206
rect 4914 2160 4920 2194
rect 4954 2160 4960 2194
rect 4914 2148 4960 2160
rect 4923 1802 4951 2148
rect 4914 1790 4960 1802
rect 4914 1756 4920 1790
rect 4954 1756 4960 1790
rect 4914 1744 4960 1756
rect 4834 1404 4880 1416
rect 4754 1217 4800 1382
rect 4834 1370 4840 1404
rect 4874 1370 4880 1404
rect 4834 1358 4880 1370
rect 4751 1211 4803 1217
rect 4751 1153 4803 1159
rect 4674 888 4720 988
rect 4674 854 4680 888
rect 4714 854 4720 888
rect 4674 822 4720 854
rect 4671 816 4723 822
rect 4671 758 4723 764
rect 4594 726 4640 738
rect 4594 692 4600 726
rect 4634 692 4640 726
rect 4594 680 4640 692
rect 4603 592 4631 680
rect 4594 427 4640 592
rect 4591 421 4643 427
rect 4591 363 4643 369
rect 1348 187 1406 193
rect 1348 153 1360 187
rect 1394 153 1406 187
rect 1348 147 1406 153
rect 4411 94 4417 146
rect 4469 94 4475 146
rect 4514 98 4560 198
rect 4514 64 4520 98
rect 4554 64 4560 98
rect 4514 32 4560 64
rect 4511 26 4563 32
rect 4603 0 4631 363
rect 4683 0 4711 758
rect 4763 0 4791 1153
rect 4843 1012 4871 1358
rect 4834 1000 4880 1012
rect 4834 966 4840 1000
rect 4874 966 4880 1000
rect 4834 954 4880 966
rect 4843 626 4871 954
rect 4834 614 4880 626
rect 4834 580 4840 614
rect 4874 580 4880 614
rect 4834 568 4880 580
rect 4843 222 4871 568
rect 4834 210 4880 222
rect 4834 176 4840 210
rect 4874 176 4880 210
rect 4834 164 4880 176
rect 4843 0 4871 164
rect 4923 0 4951 1744
rect 5003 0 5031 3128
rect 5083 0 5111 3523
rect 5163 3472 5191 3638
rect 5154 3460 5200 3472
rect 5154 3426 5160 3460
rect 5194 3426 5200 3460
rect 5154 3414 5200 3426
rect 5163 2906 5191 3414
rect 5154 2894 5200 2906
rect 5154 2860 5160 2894
rect 5194 2860 5200 2894
rect 5154 2848 5200 2860
rect 5163 2682 5191 2848
rect 5154 2670 5200 2682
rect 5154 2636 5160 2670
rect 5194 2636 5200 2670
rect 5154 2624 5200 2636
rect 5163 2116 5191 2624
rect 5154 2104 5200 2116
rect 5154 2070 5160 2104
rect 5194 2070 5200 2104
rect 5154 2058 5200 2070
rect 5163 1892 5191 2058
rect 5154 1880 5200 1892
rect 5154 1846 5160 1880
rect 5194 1846 5200 1880
rect 5154 1834 5200 1846
rect 5163 1326 5191 1834
rect 5154 1314 5200 1326
rect 5154 1280 5160 1314
rect 5194 1280 5200 1314
rect 5154 1268 5200 1280
rect 5163 1102 5191 1268
rect 5154 1090 5200 1102
rect 5154 1056 5160 1090
rect 5194 1056 5200 1090
rect 5154 1044 5200 1056
rect 5163 536 5191 1044
rect 5154 524 5200 536
rect 5154 490 5160 524
rect 5194 490 5200 524
rect 5154 478 5200 490
rect 5163 312 5191 478
rect 5154 300 5200 312
rect 5154 266 5160 300
rect 5194 266 5200 300
rect 5154 254 5200 266
rect 5163 0 5191 254
rect 5243 0 5271 5103
rect 5323 0 5351 5498
rect 5403 0 5431 5893
rect 5483 0 5511 6288
rect 5563 0 5591 6683
rect 5643 0 5671 7078
rect 5723 0 5751 7473
rect 6051 7180 6097 7502
rect 6042 7128 6048 7180
rect 6100 7128 6106 7180
rect 6051 6764 6097 7128
rect 6475 7122 6523 7502
rect 6907 7122 6955 7502
rect 7281 7479 7287 7531
rect 7339 7479 7345 7531
rect 7677 7479 7683 7531
rect 7735 7479 7741 7531
rect 7299 7136 7327 7479
rect 7695 7136 7723 7479
rect 6467 7070 6473 7122
rect 6525 7070 6531 7122
rect 6899 7070 6905 7122
rect 6957 7070 6963 7122
rect 7281 7084 7287 7136
rect 7339 7084 7345 7136
rect 7677 7084 7683 7136
rect 7735 7084 7741 7136
rect 6475 6764 6523 7070
rect 6907 6764 6955 7070
rect 6042 6712 6048 6764
rect 6100 6712 6106 6764
rect 6467 6712 6473 6764
rect 6525 6712 6531 6764
rect 6899 6712 6905 6764
rect 6957 6712 6963 6764
rect 7299 6741 7327 7084
rect 7695 6741 7723 7084
rect 6051 6390 6097 6712
rect 6042 6338 6048 6390
rect 6100 6338 6106 6390
rect 6051 5974 6097 6338
rect 6475 6332 6523 6712
rect 6907 6332 6955 6712
rect 7281 6689 7287 6741
rect 7339 6689 7345 6741
rect 7677 6689 7683 6741
rect 7735 6689 7741 6741
rect 7299 6346 7327 6689
rect 7695 6346 7723 6689
rect 6467 6280 6473 6332
rect 6525 6280 6531 6332
rect 6899 6280 6905 6332
rect 6957 6280 6963 6332
rect 7281 6294 7287 6346
rect 7339 6294 7345 6346
rect 7677 6294 7683 6346
rect 7735 6294 7741 6346
rect 6475 5974 6523 6280
rect 6907 5974 6955 6280
rect 6042 5922 6048 5974
rect 6100 5922 6106 5974
rect 6467 5922 6473 5974
rect 6525 5922 6531 5974
rect 6899 5922 6905 5974
rect 6957 5922 6963 5974
rect 7299 5951 7327 6294
rect 7695 5951 7723 6294
rect 6051 5600 6097 5922
rect 6042 5548 6048 5600
rect 6100 5548 6106 5600
rect 6051 5184 6097 5548
rect 6475 5542 6523 5922
rect 6907 5542 6955 5922
rect 7281 5899 7287 5951
rect 7339 5899 7345 5951
rect 7677 5899 7683 5951
rect 7735 5899 7741 5951
rect 7299 5556 7327 5899
rect 7695 5556 7723 5899
rect 6467 5490 6473 5542
rect 6525 5490 6531 5542
rect 6899 5490 6905 5542
rect 6957 5490 6963 5542
rect 7281 5504 7287 5556
rect 7339 5504 7345 5556
rect 7677 5504 7683 5556
rect 7735 5504 7741 5556
rect 6475 5184 6523 5490
rect 6907 5184 6955 5490
rect 6042 5132 6048 5184
rect 6100 5132 6106 5184
rect 6467 5132 6473 5184
rect 6525 5132 6531 5184
rect 6899 5132 6905 5184
rect 6957 5132 6963 5184
rect 7299 5161 7327 5504
rect 7695 5161 7723 5504
rect 6051 4810 6097 5132
rect 6042 4758 6048 4810
rect 6100 4758 6106 4810
rect 6051 4394 6097 4758
rect 6475 4752 6523 5132
rect 6907 4752 6955 5132
rect 7281 5109 7287 5161
rect 7339 5109 7345 5161
rect 7677 5109 7683 5161
rect 7735 5109 7741 5161
rect 7299 4766 7327 5109
rect 7695 4766 7723 5109
rect 6467 4700 6473 4752
rect 6525 4700 6531 4752
rect 6899 4700 6905 4752
rect 6957 4700 6963 4752
rect 7281 4714 7287 4766
rect 7339 4714 7345 4766
rect 7677 4714 7683 4766
rect 7735 4714 7741 4766
rect 6475 4394 6523 4700
rect 6907 4394 6955 4700
rect 6042 4342 6048 4394
rect 6100 4342 6106 4394
rect 6467 4342 6473 4394
rect 6525 4342 6531 4394
rect 6899 4342 6905 4394
rect 6957 4342 6963 4394
rect 7299 4371 7327 4714
rect 7695 4371 7723 4714
rect 6051 4020 6097 4342
rect 6042 3968 6048 4020
rect 6100 3968 6106 4020
rect 6051 3604 6097 3968
rect 6475 3962 6523 4342
rect 6907 3962 6955 4342
rect 7281 4319 7287 4371
rect 7339 4319 7345 4371
rect 7677 4319 7683 4371
rect 7735 4319 7741 4371
rect 7299 3976 7327 4319
rect 7695 3976 7723 4319
rect 6467 3910 6473 3962
rect 6525 3910 6531 3962
rect 6899 3910 6905 3962
rect 6957 3910 6963 3962
rect 7281 3924 7287 3976
rect 7339 3924 7345 3976
rect 7677 3924 7683 3976
rect 7735 3924 7741 3976
rect 6475 3604 6523 3910
rect 6907 3604 6955 3910
rect 6042 3552 6048 3604
rect 6100 3552 6106 3604
rect 6467 3552 6473 3604
rect 6525 3552 6531 3604
rect 6899 3552 6905 3604
rect 6957 3552 6963 3604
rect 7299 3581 7327 3924
rect 7695 3581 7723 3924
rect 6051 3230 6097 3552
rect 6042 3178 6048 3230
rect 6100 3178 6106 3230
rect 6051 2814 6097 3178
rect 6475 3172 6523 3552
rect 6907 3172 6955 3552
rect 7281 3529 7287 3581
rect 7339 3529 7345 3581
rect 7677 3529 7683 3581
rect 7735 3529 7741 3581
rect 7299 3186 7327 3529
rect 7695 3186 7723 3529
rect 6467 3120 6473 3172
rect 6525 3120 6531 3172
rect 6899 3120 6905 3172
rect 6957 3120 6963 3172
rect 7281 3134 7287 3186
rect 7339 3134 7345 3186
rect 7677 3134 7683 3186
rect 7735 3134 7741 3186
rect 6475 2814 6523 3120
rect 6907 2814 6955 3120
rect 6042 2762 6048 2814
rect 6100 2762 6106 2814
rect 6467 2762 6473 2814
rect 6525 2762 6531 2814
rect 6899 2762 6905 2814
rect 6957 2762 6963 2814
rect 7299 2791 7327 3134
rect 7695 2791 7723 3134
rect 6051 2440 6097 2762
rect 6042 2388 6048 2440
rect 6100 2388 6106 2440
rect 6051 2024 6097 2388
rect 6475 2382 6523 2762
rect 6907 2382 6955 2762
rect 7281 2739 7287 2791
rect 7339 2739 7345 2791
rect 7677 2739 7683 2791
rect 7735 2739 7741 2791
rect 7299 2396 7327 2739
rect 7695 2396 7723 2739
rect 6467 2330 6473 2382
rect 6525 2330 6531 2382
rect 6899 2330 6905 2382
rect 6957 2330 6963 2382
rect 7281 2344 7287 2396
rect 7339 2344 7345 2396
rect 7677 2344 7683 2396
rect 7735 2344 7741 2396
rect 6475 2024 6523 2330
rect 6907 2024 6955 2330
rect 6042 1972 6048 2024
rect 6100 1972 6106 2024
rect 6467 1972 6473 2024
rect 6525 1972 6531 2024
rect 6899 1972 6905 2024
rect 6957 1972 6963 2024
rect 7299 2001 7327 2344
rect 7695 2001 7723 2344
rect 6051 1650 6097 1972
rect 6042 1598 6048 1650
rect 6100 1598 6106 1650
rect 6051 1234 6097 1598
rect 6475 1592 6523 1972
rect 6907 1592 6955 1972
rect 7281 1949 7287 2001
rect 7339 1949 7345 2001
rect 7677 1949 7683 2001
rect 7735 1949 7741 2001
rect 7299 1606 7327 1949
rect 7695 1606 7723 1949
rect 6467 1540 6473 1592
rect 6525 1540 6531 1592
rect 6899 1540 6905 1592
rect 6957 1540 6963 1592
rect 7281 1554 7287 1606
rect 7339 1554 7345 1606
rect 7677 1554 7683 1606
rect 7735 1554 7741 1606
rect 6475 1234 6523 1540
rect 6907 1234 6955 1540
rect 6042 1182 6048 1234
rect 6100 1182 6106 1234
rect 6467 1182 6473 1234
rect 6525 1182 6531 1234
rect 6899 1182 6905 1234
rect 6957 1182 6963 1234
rect 7299 1211 7327 1554
rect 7695 1211 7723 1554
rect 6051 860 6097 1182
rect 6042 808 6048 860
rect 6100 808 6106 860
rect 6051 444 6097 808
rect 6475 802 6523 1182
rect 6907 802 6955 1182
rect 7281 1159 7287 1211
rect 7339 1159 7345 1211
rect 7677 1159 7683 1211
rect 7735 1159 7741 1211
rect 7299 816 7327 1159
rect 7695 816 7723 1159
rect 6467 750 6473 802
rect 6525 750 6531 802
rect 6899 750 6905 802
rect 6957 750 6963 802
rect 7281 764 7287 816
rect 7339 764 7345 816
rect 7677 764 7683 816
rect 7735 764 7741 816
rect 6475 444 6523 750
rect 6907 444 6955 750
rect 6042 392 6048 444
rect 6100 392 6106 444
rect 6467 392 6473 444
rect 6525 392 6531 444
rect 6899 392 6905 444
rect 6957 392 6963 444
rect 7299 421 7327 764
rect 7695 421 7723 764
rect 6051 -16 6097 392
rect 6475 42 6523 392
rect 6907 42 6955 392
rect 7281 369 7287 421
rect 7339 369 7345 421
rect 7677 369 7683 421
rect 7735 369 7741 421
rect 7299 28 7327 369
rect 7695 28 7723 369
rect 4511 -32 4563 -26
<< via1 >>
rect 4417 7797 4469 7806
rect 4417 7763 4426 7797
rect 4426 7763 4460 7797
rect 4460 7763 4469 7797
rect 4417 7754 4469 7763
rect 4417 7247 4469 7256
rect 4417 7213 4426 7247
rect 4426 7213 4460 7247
rect 4460 7213 4469 7247
rect 4417 7204 4469 7213
rect 4417 7007 4469 7016
rect 4417 6973 4426 7007
rect 4426 6973 4460 7007
rect 4460 6973 4469 7007
rect 4417 6964 4469 6973
rect 4417 6457 4469 6466
rect 4417 6423 4426 6457
rect 4426 6423 4460 6457
rect 4460 6423 4469 6457
rect 4417 6414 4469 6423
rect 4417 6217 4469 6226
rect 4417 6183 4426 6217
rect 4426 6183 4460 6217
rect 4460 6183 4469 6217
rect 4417 6174 4469 6183
rect 4417 5667 4469 5676
rect 4417 5633 4426 5667
rect 4426 5633 4460 5667
rect 4460 5633 4469 5667
rect 4417 5624 4469 5633
rect 4417 5427 4469 5436
rect 4417 5393 4426 5427
rect 4426 5393 4460 5427
rect 4460 5393 4469 5427
rect 4417 5384 4469 5393
rect 4417 4877 4469 4886
rect 4417 4843 4426 4877
rect 4426 4843 4460 4877
rect 4460 4843 4469 4877
rect 4417 4834 4469 4843
rect 4417 3847 4469 3856
rect 4417 3813 4426 3847
rect 4426 3813 4460 3847
rect 4460 3813 4469 3847
rect 4417 3804 4469 3813
rect 4417 3297 4469 3306
rect 4417 3263 4426 3297
rect 4426 3263 4460 3297
rect 4460 3263 4469 3297
rect 4417 3254 4469 3263
rect 4417 3057 4469 3066
rect 4417 3023 4426 3057
rect 4426 3023 4460 3057
rect 4460 3023 4469 3057
rect 4417 3014 4469 3023
rect 4417 2507 4469 2516
rect 4417 2473 4426 2507
rect 4426 2473 4460 2507
rect 4460 2473 4469 2507
rect 4417 2464 4469 2473
rect 4417 1477 4469 1486
rect 4417 1443 4426 1477
rect 4426 1443 4460 1477
rect 4460 1443 4469 1477
rect 4417 1434 4469 1443
rect 4417 927 4469 936
rect 4417 893 4426 927
rect 4426 893 4460 927
rect 4460 893 4469 927
rect 4417 884 4469 893
rect 4417 687 4469 696
rect 4417 653 4426 687
rect 4426 653 4460 687
rect 4460 653 4469 687
rect 4417 644 4469 653
rect 6048 50162 6100 50214
rect 6473 50162 6525 50214
rect 6905 50162 6957 50214
rect 6048 49788 6100 49840
rect 7287 50139 7339 50191
rect 7683 50139 7735 50191
rect 6473 49730 6525 49782
rect 6905 49730 6957 49782
rect 7287 49744 7339 49796
rect 7683 49744 7735 49796
rect 6048 49372 6100 49424
rect 6473 49372 6525 49424
rect 6905 49372 6957 49424
rect 6048 48998 6100 49050
rect 7287 49349 7339 49401
rect 7683 49349 7735 49401
rect 6473 48940 6525 48992
rect 6905 48940 6957 48992
rect 7287 48954 7339 49006
rect 7683 48954 7735 49006
rect 6048 48582 6100 48634
rect 6473 48582 6525 48634
rect 6905 48582 6957 48634
rect 6048 48208 6100 48260
rect 7287 48559 7339 48611
rect 7683 48559 7735 48611
rect 6473 48150 6525 48202
rect 6905 48150 6957 48202
rect 7287 48164 7339 48216
rect 7683 48164 7735 48216
rect 6048 47792 6100 47844
rect 6473 47792 6525 47844
rect 6905 47792 6957 47844
rect 6048 47418 6100 47470
rect 7287 47769 7339 47821
rect 7683 47769 7735 47821
rect 6473 47360 6525 47412
rect 6905 47360 6957 47412
rect 7287 47374 7339 47426
rect 7683 47374 7735 47426
rect 6048 47002 6100 47054
rect 6473 47002 6525 47054
rect 6905 47002 6957 47054
rect 6048 46628 6100 46680
rect 7287 46979 7339 47031
rect 7683 46979 7735 47031
rect 6473 46570 6525 46622
rect 6905 46570 6957 46622
rect 7287 46584 7339 46636
rect 7683 46584 7735 46636
rect 6048 46212 6100 46264
rect 6473 46212 6525 46264
rect 6905 46212 6957 46264
rect 6048 45838 6100 45890
rect 7287 46189 7339 46241
rect 7683 46189 7735 46241
rect 6473 45780 6525 45832
rect 6905 45780 6957 45832
rect 7287 45794 7339 45846
rect 7683 45794 7735 45846
rect 6048 45422 6100 45474
rect 6473 45422 6525 45474
rect 6905 45422 6957 45474
rect 6048 45048 6100 45100
rect 7287 45399 7339 45451
rect 7683 45399 7735 45451
rect 6473 44990 6525 45042
rect 6905 44990 6957 45042
rect 7287 45004 7339 45056
rect 7683 45004 7735 45056
rect 6048 44632 6100 44684
rect 6473 44632 6525 44684
rect 6905 44632 6957 44684
rect 6048 44258 6100 44310
rect 7287 44609 7339 44661
rect 7683 44609 7735 44661
rect 6473 44200 6525 44252
rect 6905 44200 6957 44252
rect 7287 44214 7339 44266
rect 7683 44214 7735 44266
rect 6048 43842 6100 43894
rect 6473 43842 6525 43894
rect 6905 43842 6957 43894
rect 6048 43468 6100 43520
rect 7287 43819 7339 43871
rect 7683 43819 7735 43871
rect 6473 43410 6525 43462
rect 6905 43410 6957 43462
rect 7287 43424 7339 43476
rect 7683 43424 7735 43476
rect 6048 43052 6100 43104
rect 6473 43052 6525 43104
rect 6905 43052 6957 43104
rect 6048 42678 6100 42730
rect 7287 43029 7339 43081
rect 7683 43029 7735 43081
rect 6473 42620 6525 42672
rect 6905 42620 6957 42672
rect 7287 42634 7339 42686
rect 7683 42634 7735 42686
rect 6048 42262 6100 42314
rect 6473 42262 6525 42314
rect 6905 42262 6957 42314
rect 6048 41888 6100 41940
rect 7287 42239 7339 42291
rect 7683 42239 7735 42291
rect 6473 41830 6525 41882
rect 6905 41830 6957 41882
rect 7287 41844 7339 41896
rect 7683 41844 7735 41896
rect 6048 41472 6100 41524
rect 6473 41472 6525 41524
rect 6905 41472 6957 41524
rect 6048 41098 6100 41150
rect 7287 41449 7339 41501
rect 7683 41449 7735 41501
rect 6473 41040 6525 41092
rect 6905 41040 6957 41092
rect 7287 41054 7339 41106
rect 7683 41054 7735 41106
rect 6048 40682 6100 40734
rect 6473 40682 6525 40734
rect 6905 40682 6957 40734
rect 6048 40308 6100 40360
rect 7287 40659 7339 40711
rect 7683 40659 7735 40711
rect 6473 40250 6525 40302
rect 6905 40250 6957 40302
rect 7287 40264 7339 40316
rect 7683 40264 7735 40316
rect 6048 39892 6100 39944
rect 6473 39892 6525 39944
rect 6905 39892 6957 39944
rect 6048 39518 6100 39570
rect 7287 39869 7339 39921
rect 7683 39869 7735 39921
rect 6473 39460 6525 39512
rect 6905 39460 6957 39512
rect 7287 39474 7339 39526
rect 7683 39474 7735 39526
rect 6048 39102 6100 39154
rect 6473 39102 6525 39154
rect 6905 39102 6957 39154
rect 6048 38728 6100 38780
rect 7287 39079 7339 39131
rect 7683 39079 7735 39131
rect 6473 38670 6525 38722
rect 6905 38670 6957 38722
rect 7287 38684 7339 38736
rect 7683 38684 7735 38736
rect 6048 38312 6100 38364
rect 6473 38312 6525 38364
rect 6905 38312 6957 38364
rect 6048 37938 6100 37990
rect 7287 38289 7339 38341
rect 7683 38289 7735 38341
rect 6473 37880 6525 37932
rect 6905 37880 6957 37932
rect 7287 37894 7339 37946
rect 7683 37894 7735 37946
rect 6048 37522 6100 37574
rect 6473 37522 6525 37574
rect 6905 37522 6957 37574
rect 6048 37148 6100 37200
rect 7287 37499 7339 37551
rect 7683 37499 7735 37551
rect 6473 37090 6525 37142
rect 6905 37090 6957 37142
rect 7287 37104 7339 37156
rect 7683 37104 7735 37156
rect 6048 36732 6100 36784
rect 6473 36732 6525 36784
rect 6905 36732 6957 36784
rect 6048 36358 6100 36410
rect 7287 36709 7339 36761
rect 7683 36709 7735 36761
rect 6473 36300 6525 36352
rect 6905 36300 6957 36352
rect 7287 36314 7339 36366
rect 7683 36314 7735 36366
rect 6048 35942 6100 35994
rect 6473 35942 6525 35994
rect 6905 35942 6957 35994
rect 6048 35568 6100 35620
rect 7287 35919 7339 35971
rect 7683 35919 7735 35971
rect 6473 35510 6525 35562
rect 6905 35510 6957 35562
rect 7287 35524 7339 35576
rect 7683 35524 7735 35576
rect 6048 35152 6100 35204
rect 6473 35152 6525 35204
rect 6905 35152 6957 35204
rect 6048 34778 6100 34830
rect 7287 35129 7339 35181
rect 7683 35129 7735 35181
rect 6473 34720 6525 34772
rect 6905 34720 6957 34772
rect 7287 34734 7339 34786
rect 7683 34734 7735 34786
rect 6048 34362 6100 34414
rect 6473 34362 6525 34414
rect 6905 34362 6957 34414
rect 6048 33988 6100 34040
rect 7287 34339 7339 34391
rect 7683 34339 7735 34391
rect 6473 33930 6525 33982
rect 6905 33930 6957 33982
rect 7287 33944 7339 33996
rect 7683 33944 7735 33996
rect 6048 33572 6100 33624
rect 6473 33572 6525 33624
rect 6905 33572 6957 33624
rect 6048 33198 6100 33250
rect 7287 33549 7339 33601
rect 7683 33549 7735 33601
rect 6473 33140 6525 33192
rect 6905 33140 6957 33192
rect 7287 33154 7339 33206
rect 7683 33154 7735 33206
rect 6048 32782 6100 32834
rect 6473 32782 6525 32834
rect 6905 32782 6957 32834
rect 6048 32408 6100 32460
rect 7287 32759 7339 32811
rect 7683 32759 7735 32811
rect 6473 32350 6525 32402
rect 6905 32350 6957 32402
rect 7287 32364 7339 32416
rect 7683 32364 7735 32416
rect 6048 31992 6100 32044
rect 6473 31992 6525 32044
rect 6905 31992 6957 32044
rect 6048 31618 6100 31670
rect 7287 31969 7339 32021
rect 7683 31969 7735 32021
rect 6473 31560 6525 31612
rect 6905 31560 6957 31612
rect 7287 31574 7339 31626
rect 7683 31574 7735 31626
rect 6048 31202 6100 31254
rect 6473 31202 6525 31254
rect 6905 31202 6957 31254
rect 6048 30828 6100 30880
rect 7287 31179 7339 31231
rect 7683 31179 7735 31231
rect 6473 30770 6525 30822
rect 6905 30770 6957 30822
rect 7287 30784 7339 30836
rect 7683 30784 7735 30836
rect 6048 30412 6100 30464
rect 6473 30412 6525 30464
rect 6905 30412 6957 30464
rect 6048 30038 6100 30090
rect 7287 30389 7339 30441
rect 7683 30389 7735 30441
rect 6473 29980 6525 30032
rect 6905 29980 6957 30032
rect 7287 29994 7339 30046
rect 7683 29994 7735 30046
rect 6048 29622 6100 29674
rect 6473 29622 6525 29674
rect 6905 29622 6957 29674
rect 6048 29248 6100 29300
rect 7287 29599 7339 29651
rect 7683 29599 7735 29651
rect 6473 29190 6525 29242
rect 6905 29190 6957 29242
rect 7287 29204 7339 29256
rect 7683 29204 7735 29256
rect 6048 28832 6100 28884
rect 6473 28832 6525 28884
rect 6905 28832 6957 28884
rect 6048 28458 6100 28510
rect 7287 28809 7339 28861
rect 7683 28809 7735 28861
rect 6473 28400 6525 28452
rect 6905 28400 6957 28452
rect 7287 28414 7339 28466
rect 7683 28414 7735 28466
rect 6048 28042 6100 28094
rect 6473 28042 6525 28094
rect 6905 28042 6957 28094
rect 6048 27668 6100 27720
rect 7287 28019 7339 28071
rect 7683 28019 7735 28071
rect 6473 27610 6525 27662
rect 6905 27610 6957 27662
rect 7287 27624 7339 27676
rect 7683 27624 7735 27676
rect 6048 27252 6100 27304
rect 6473 27252 6525 27304
rect 6905 27252 6957 27304
rect 6048 26878 6100 26930
rect 7287 27229 7339 27281
rect 7683 27229 7735 27281
rect 6473 26820 6525 26872
rect 6905 26820 6957 26872
rect 7287 26834 7339 26886
rect 7683 26834 7735 26886
rect 6048 26462 6100 26514
rect 6473 26462 6525 26514
rect 6905 26462 6957 26514
rect 6048 26088 6100 26140
rect 7287 26439 7339 26491
rect 7683 26439 7735 26491
rect 6473 26030 6525 26082
rect 6905 26030 6957 26082
rect 7287 26044 7339 26096
rect 7683 26044 7735 26096
rect 6048 25672 6100 25724
rect 6473 25672 6525 25724
rect 6905 25672 6957 25724
rect 6048 25298 6100 25350
rect 7287 25649 7339 25701
rect 7683 25649 7735 25701
rect 6473 25240 6525 25292
rect 6905 25240 6957 25292
rect 7287 25254 7339 25306
rect 7683 25254 7735 25306
rect 6048 24882 6100 24934
rect 6473 24882 6525 24934
rect 6905 24882 6957 24934
rect 6048 24508 6100 24560
rect 7287 24859 7339 24911
rect 7683 24859 7735 24911
rect 6473 24450 6525 24502
rect 6905 24450 6957 24502
rect 7287 24464 7339 24516
rect 7683 24464 7735 24516
rect 6048 24092 6100 24144
rect 6473 24092 6525 24144
rect 6905 24092 6957 24144
rect 6048 23718 6100 23770
rect 7287 24069 7339 24121
rect 7683 24069 7735 24121
rect 6473 23660 6525 23712
rect 6905 23660 6957 23712
rect 7287 23674 7339 23726
rect 7683 23674 7735 23726
rect 6048 23302 6100 23354
rect 6473 23302 6525 23354
rect 6905 23302 6957 23354
rect 6048 22928 6100 22980
rect 7287 23279 7339 23331
rect 7683 23279 7735 23331
rect 6473 22870 6525 22922
rect 6905 22870 6957 22922
rect 7287 22884 7339 22936
rect 7683 22884 7735 22936
rect 6048 22512 6100 22564
rect 6473 22512 6525 22564
rect 6905 22512 6957 22564
rect 6048 22138 6100 22190
rect 7287 22489 7339 22541
rect 7683 22489 7735 22541
rect 6473 22080 6525 22132
rect 6905 22080 6957 22132
rect 7287 22094 7339 22146
rect 7683 22094 7735 22146
rect 6048 21722 6100 21774
rect 6473 21722 6525 21774
rect 6905 21722 6957 21774
rect 6048 21348 6100 21400
rect 7287 21699 7339 21751
rect 7683 21699 7735 21751
rect 6473 21290 6525 21342
rect 6905 21290 6957 21342
rect 7287 21304 7339 21356
rect 7683 21304 7735 21356
rect 6048 20932 6100 20984
rect 6473 20932 6525 20984
rect 6905 20932 6957 20984
rect 6048 20558 6100 20610
rect 7287 20909 7339 20961
rect 7683 20909 7735 20961
rect 6473 20500 6525 20552
rect 6905 20500 6957 20552
rect 7287 20514 7339 20566
rect 7683 20514 7735 20566
rect 6048 20142 6100 20194
rect 6473 20142 6525 20194
rect 6905 20142 6957 20194
rect 6048 19768 6100 19820
rect 7287 20119 7339 20171
rect 7683 20119 7735 20171
rect 6473 19710 6525 19762
rect 6905 19710 6957 19762
rect 7287 19724 7339 19776
rect 7683 19724 7735 19776
rect 6048 19352 6100 19404
rect 6473 19352 6525 19404
rect 6905 19352 6957 19404
rect 6048 18978 6100 19030
rect 7287 19329 7339 19381
rect 7683 19329 7735 19381
rect 6473 18920 6525 18972
rect 6905 18920 6957 18972
rect 7287 18934 7339 18986
rect 7683 18934 7735 18986
rect 6048 18562 6100 18614
rect 6473 18562 6525 18614
rect 6905 18562 6957 18614
rect 6048 18188 6100 18240
rect 7287 18539 7339 18591
rect 7683 18539 7735 18591
rect 6473 18130 6525 18182
rect 6905 18130 6957 18182
rect 7287 18144 7339 18196
rect 7683 18144 7735 18196
rect 6048 17772 6100 17824
rect 6473 17772 6525 17824
rect 6905 17772 6957 17824
rect 6048 17398 6100 17450
rect 7287 17749 7339 17801
rect 7683 17749 7735 17801
rect 6473 17340 6525 17392
rect 6905 17340 6957 17392
rect 7287 17354 7339 17406
rect 7683 17354 7735 17406
rect 6048 16982 6100 17034
rect 6473 16982 6525 17034
rect 6905 16982 6957 17034
rect 6048 16608 6100 16660
rect 7287 16959 7339 17011
rect 7683 16959 7735 17011
rect 6473 16550 6525 16602
rect 6905 16550 6957 16602
rect 7287 16564 7339 16616
rect 7683 16564 7735 16616
rect 6048 16192 6100 16244
rect 6473 16192 6525 16244
rect 6905 16192 6957 16244
rect 6048 15818 6100 15870
rect 7287 16169 7339 16221
rect 7683 16169 7735 16221
rect 6473 15760 6525 15812
rect 6905 15760 6957 15812
rect 7287 15774 7339 15826
rect 7683 15774 7735 15826
rect 6048 15402 6100 15454
rect 6473 15402 6525 15454
rect 6905 15402 6957 15454
rect 6048 15028 6100 15080
rect 7287 15379 7339 15431
rect 7683 15379 7735 15431
rect 6473 14970 6525 15022
rect 6905 14970 6957 15022
rect 7287 14984 7339 15036
rect 7683 14984 7735 15036
rect 6048 14612 6100 14664
rect 6473 14612 6525 14664
rect 6905 14612 6957 14664
rect 6048 14238 6100 14290
rect 7287 14589 7339 14641
rect 7683 14589 7735 14641
rect 6473 14180 6525 14232
rect 6905 14180 6957 14232
rect 7287 14194 7339 14246
rect 7683 14194 7735 14246
rect 6048 13822 6100 13874
rect 6473 13822 6525 13874
rect 6905 13822 6957 13874
rect 6048 13448 6100 13500
rect 7287 13799 7339 13851
rect 7683 13799 7735 13851
rect 6473 13390 6525 13442
rect 6905 13390 6957 13442
rect 7287 13404 7339 13456
rect 7683 13404 7735 13456
rect 6048 13032 6100 13084
rect 6473 13032 6525 13084
rect 6905 13032 6957 13084
rect 6048 12658 6100 12710
rect 7287 13009 7339 13061
rect 7683 13009 7735 13061
rect 6473 12600 6525 12652
rect 6905 12600 6957 12652
rect 7287 12614 7339 12666
rect 7683 12614 7735 12666
rect 6048 12242 6100 12294
rect 6473 12242 6525 12294
rect 6905 12242 6957 12294
rect 6048 11868 6100 11920
rect 7287 12219 7339 12271
rect 7683 12219 7735 12271
rect 6473 11810 6525 11862
rect 6905 11810 6957 11862
rect 7287 11824 7339 11876
rect 7683 11824 7735 11876
rect 6048 11452 6100 11504
rect 6473 11452 6525 11504
rect 6905 11452 6957 11504
rect 6048 11078 6100 11130
rect 7287 11429 7339 11481
rect 7683 11429 7735 11481
rect 6473 11020 6525 11072
rect 6905 11020 6957 11072
rect 7287 11034 7339 11086
rect 7683 11034 7735 11086
rect 6048 10662 6100 10714
rect 6473 10662 6525 10714
rect 6905 10662 6957 10714
rect 6048 10288 6100 10340
rect 7287 10639 7339 10691
rect 7683 10639 7735 10691
rect 6473 10230 6525 10282
rect 6905 10230 6957 10282
rect 7287 10244 7339 10296
rect 7683 10244 7735 10296
rect 6048 9872 6100 9924
rect 6473 9872 6525 9924
rect 6905 9872 6957 9924
rect 6048 9498 6100 9550
rect 7287 9849 7339 9901
rect 7683 9849 7735 9901
rect 6473 9440 6525 9492
rect 6905 9440 6957 9492
rect 7287 9454 7339 9506
rect 7683 9454 7735 9506
rect 6048 9082 6100 9134
rect 6473 9082 6525 9134
rect 6905 9082 6957 9134
rect 6048 8708 6100 8760
rect 7287 9059 7339 9111
rect 7683 9059 7735 9111
rect 6473 8650 6525 8702
rect 6905 8650 6957 8702
rect 7287 8664 7339 8716
rect 7683 8664 7735 8716
rect 6048 8292 6100 8344
rect 6473 8292 6525 8344
rect 6905 8292 6957 8344
rect 6048 7918 6100 7970
rect 7287 8269 7339 8321
rect 7683 8269 7735 8321
rect 6473 7860 6525 7912
rect 6905 7860 6957 7912
rect 7287 7874 7339 7926
rect 7683 7874 7735 7926
rect 5711 7479 5763 7531
rect 6048 7502 6100 7554
rect 6473 7502 6525 7554
rect 6905 7502 6957 7554
rect 5631 7084 5683 7136
rect 5551 6689 5603 6741
rect 5471 6294 5523 6346
rect 5391 5899 5443 5951
rect 5311 5504 5363 5556
rect 5231 5109 5283 5161
rect 5151 4714 5203 4766
rect 5071 3529 5123 3581
rect 4991 3134 5043 3186
rect 4911 2739 4963 2791
rect 4831 2344 4883 2396
rect 4751 1159 4803 1211
rect 4671 764 4723 816
rect 4591 369 4643 421
rect 4417 137 4469 146
rect 4417 103 4426 137
rect 4426 103 4460 137
rect 4460 103 4469 137
rect 4417 94 4469 103
rect 4511 -26 4563 26
rect 6048 7128 6100 7180
rect 7287 7479 7339 7531
rect 7683 7479 7735 7531
rect 6473 7070 6525 7122
rect 6905 7070 6957 7122
rect 7287 7084 7339 7136
rect 7683 7084 7735 7136
rect 6048 6712 6100 6764
rect 6473 6712 6525 6764
rect 6905 6712 6957 6764
rect 6048 6338 6100 6390
rect 7287 6689 7339 6741
rect 7683 6689 7735 6741
rect 6473 6280 6525 6332
rect 6905 6280 6957 6332
rect 7287 6294 7339 6346
rect 7683 6294 7735 6346
rect 6048 5922 6100 5974
rect 6473 5922 6525 5974
rect 6905 5922 6957 5974
rect 6048 5548 6100 5600
rect 7287 5899 7339 5951
rect 7683 5899 7735 5951
rect 6473 5490 6525 5542
rect 6905 5490 6957 5542
rect 7287 5504 7339 5556
rect 7683 5504 7735 5556
rect 6048 5132 6100 5184
rect 6473 5132 6525 5184
rect 6905 5132 6957 5184
rect 6048 4758 6100 4810
rect 7287 5109 7339 5161
rect 7683 5109 7735 5161
rect 6473 4700 6525 4752
rect 6905 4700 6957 4752
rect 7287 4714 7339 4766
rect 7683 4714 7735 4766
rect 6048 4342 6100 4394
rect 6473 4342 6525 4394
rect 6905 4342 6957 4394
rect 6048 3968 6100 4020
rect 7287 4319 7339 4371
rect 7683 4319 7735 4371
rect 6473 3910 6525 3962
rect 6905 3910 6957 3962
rect 7287 3924 7339 3976
rect 7683 3924 7735 3976
rect 6048 3552 6100 3604
rect 6473 3552 6525 3604
rect 6905 3552 6957 3604
rect 6048 3178 6100 3230
rect 7287 3529 7339 3581
rect 7683 3529 7735 3581
rect 6473 3120 6525 3172
rect 6905 3120 6957 3172
rect 7287 3134 7339 3186
rect 7683 3134 7735 3186
rect 6048 2762 6100 2814
rect 6473 2762 6525 2814
rect 6905 2762 6957 2814
rect 6048 2388 6100 2440
rect 7287 2739 7339 2791
rect 7683 2739 7735 2791
rect 6473 2330 6525 2382
rect 6905 2330 6957 2382
rect 7287 2344 7339 2396
rect 7683 2344 7735 2396
rect 6048 1972 6100 2024
rect 6473 1972 6525 2024
rect 6905 1972 6957 2024
rect 6048 1598 6100 1650
rect 7287 1949 7339 2001
rect 7683 1949 7735 2001
rect 6473 1540 6525 1592
rect 6905 1540 6957 1592
rect 7287 1554 7339 1606
rect 7683 1554 7735 1606
rect 6048 1182 6100 1234
rect 6473 1182 6525 1234
rect 6905 1182 6957 1234
rect 6048 808 6100 860
rect 7287 1159 7339 1211
rect 7683 1159 7735 1211
rect 6473 750 6525 802
rect 6905 750 6957 802
rect 7287 764 7339 816
rect 7683 764 7735 816
rect 6048 392 6100 444
rect 6473 392 6525 444
rect 6905 392 6957 444
rect 7287 369 7339 421
rect 7683 369 7735 421
<< metal2 >>
rect 6046 50216 6102 50225
rect 6046 50151 6102 50160
rect 6471 50216 6527 50225
rect 6471 50151 6527 50160
rect 6903 50216 6959 50225
rect 6903 50151 6959 50160
rect 7285 50193 7341 50202
rect 7285 50128 7341 50137
rect 7681 50193 7737 50202
rect 7681 50128 7737 50137
rect 6046 49842 6102 49851
rect 7285 49798 7341 49807
rect 6046 49777 6102 49786
rect 6471 49784 6527 49793
rect 6471 49719 6527 49728
rect 6903 49784 6959 49793
rect 7285 49733 7341 49742
rect 7681 49798 7737 49807
rect 7681 49733 7737 49742
rect 6903 49719 6959 49728
rect 6046 49426 6102 49435
rect 6046 49361 6102 49370
rect 6471 49426 6527 49435
rect 6471 49361 6527 49370
rect 6903 49426 6959 49435
rect 6903 49361 6959 49370
rect 7285 49403 7341 49412
rect 7285 49338 7341 49347
rect 7681 49403 7737 49412
rect 7681 49338 7737 49347
rect 6046 49052 6102 49061
rect 7285 49008 7341 49017
rect 6046 48987 6102 48996
rect 6471 48994 6527 49003
rect 6471 48929 6527 48938
rect 6903 48994 6959 49003
rect 7285 48943 7341 48952
rect 7681 49008 7737 49017
rect 7681 48943 7737 48952
rect 6903 48929 6959 48938
rect 6046 48636 6102 48645
rect 6046 48571 6102 48580
rect 6471 48636 6527 48645
rect 6471 48571 6527 48580
rect 6903 48636 6959 48645
rect 6903 48571 6959 48580
rect 7285 48613 7341 48622
rect 7285 48548 7341 48557
rect 7681 48613 7737 48622
rect 7681 48548 7737 48557
rect 6046 48262 6102 48271
rect 7285 48218 7341 48227
rect 6046 48197 6102 48206
rect 6471 48204 6527 48213
rect 6471 48139 6527 48148
rect 6903 48204 6959 48213
rect 7285 48153 7341 48162
rect 7681 48218 7737 48227
rect 7681 48153 7737 48162
rect 6903 48139 6959 48148
rect 6046 47846 6102 47855
rect 6046 47781 6102 47790
rect 6471 47846 6527 47855
rect 6471 47781 6527 47790
rect 6903 47846 6959 47855
rect 6903 47781 6959 47790
rect 7285 47823 7341 47832
rect 7285 47758 7341 47767
rect 7681 47823 7737 47832
rect 7681 47758 7737 47767
rect 6046 47472 6102 47481
rect 7285 47428 7341 47437
rect 6046 47407 6102 47416
rect 6471 47414 6527 47423
rect 6471 47349 6527 47358
rect 6903 47414 6959 47423
rect 7285 47363 7341 47372
rect 7681 47428 7737 47437
rect 7681 47363 7737 47372
rect 6903 47349 6959 47358
rect 6046 47056 6102 47065
rect 6046 46991 6102 47000
rect 6471 47056 6527 47065
rect 6471 46991 6527 47000
rect 6903 47056 6959 47065
rect 6903 46991 6959 47000
rect 7285 47033 7341 47042
rect 7285 46968 7341 46977
rect 7681 47033 7737 47042
rect 7681 46968 7737 46977
rect 6046 46682 6102 46691
rect 7285 46638 7341 46647
rect 6046 46617 6102 46626
rect 6471 46624 6527 46633
rect 6471 46559 6527 46568
rect 6903 46624 6959 46633
rect 7285 46573 7341 46582
rect 7681 46638 7737 46647
rect 7681 46573 7737 46582
rect 6903 46559 6959 46568
rect 6046 46266 6102 46275
rect 6046 46201 6102 46210
rect 6471 46266 6527 46275
rect 6471 46201 6527 46210
rect 6903 46266 6959 46275
rect 6903 46201 6959 46210
rect 7285 46243 7341 46252
rect 7285 46178 7341 46187
rect 7681 46243 7737 46252
rect 7681 46178 7737 46187
rect 6046 45892 6102 45901
rect 7285 45848 7341 45857
rect 6046 45827 6102 45836
rect 6471 45834 6527 45843
rect 6471 45769 6527 45778
rect 6903 45834 6959 45843
rect 7285 45783 7341 45792
rect 7681 45848 7737 45857
rect 7681 45783 7737 45792
rect 6903 45769 6959 45778
rect 6046 45476 6102 45485
rect 6046 45411 6102 45420
rect 6471 45476 6527 45485
rect 6471 45411 6527 45420
rect 6903 45476 6959 45485
rect 6903 45411 6959 45420
rect 7285 45453 7341 45462
rect 7285 45388 7341 45397
rect 7681 45453 7737 45462
rect 7681 45388 7737 45397
rect 6046 45102 6102 45111
rect 7285 45058 7341 45067
rect 6046 45037 6102 45046
rect 6471 45044 6527 45053
rect 6471 44979 6527 44988
rect 6903 45044 6959 45053
rect 7285 44993 7341 45002
rect 7681 45058 7737 45067
rect 7681 44993 7737 45002
rect 6903 44979 6959 44988
rect 6046 44686 6102 44695
rect 6046 44621 6102 44630
rect 6471 44686 6527 44695
rect 6471 44621 6527 44630
rect 6903 44686 6959 44695
rect 6903 44621 6959 44630
rect 7285 44663 7341 44672
rect 7285 44598 7341 44607
rect 7681 44663 7737 44672
rect 7681 44598 7737 44607
rect 6046 44312 6102 44321
rect 7285 44268 7341 44277
rect 6046 44247 6102 44256
rect 6471 44254 6527 44263
rect 6471 44189 6527 44198
rect 6903 44254 6959 44263
rect 7285 44203 7341 44212
rect 7681 44268 7737 44277
rect 7681 44203 7737 44212
rect 6903 44189 6959 44198
rect 6046 43896 6102 43905
rect 6046 43831 6102 43840
rect 6471 43896 6527 43905
rect 6471 43831 6527 43840
rect 6903 43896 6959 43905
rect 6903 43831 6959 43840
rect 7285 43873 7341 43882
rect 7285 43808 7341 43817
rect 7681 43873 7737 43882
rect 7681 43808 7737 43817
rect 6046 43522 6102 43531
rect 7285 43478 7341 43487
rect 6046 43457 6102 43466
rect 6471 43464 6527 43473
rect 6471 43399 6527 43408
rect 6903 43464 6959 43473
rect 7285 43413 7341 43422
rect 7681 43478 7737 43487
rect 7681 43413 7737 43422
rect 6903 43399 6959 43408
rect 6046 43106 6102 43115
rect 6046 43041 6102 43050
rect 6471 43106 6527 43115
rect 6471 43041 6527 43050
rect 6903 43106 6959 43115
rect 6903 43041 6959 43050
rect 7285 43083 7341 43092
rect 7285 43018 7341 43027
rect 7681 43083 7737 43092
rect 7681 43018 7737 43027
rect 6046 42732 6102 42741
rect 7285 42688 7341 42697
rect 6046 42667 6102 42676
rect 6471 42674 6527 42683
rect 6471 42609 6527 42618
rect 6903 42674 6959 42683
rect 7285 42623 7341 42632
rect 7681 42688 7737 42697
rect 7681 42623 7737 42632
rect 6903 42609 6959 42618
rect 6046 42316 6102 42325
rect 6046 42251 6102 42260
rect 6471 42316 6527 42325
rect 6471 42251 6527 42260
rect 6903 42316 6959 42325
rect 6903 42251 6959 42260
rect 7285 42293 7341 42302
rect 7285 42228 7341 42237
rect 7681 42293 7737 42302
rect 7681 42228 7737 42237
rect 6046 41942 6102 41951
rect 7285 41898 7341 41907
rect 6046 41877 6102 41886
rect 6471 41884 6527 41893
rect 6471 41819 6527 41828
rect 6903 41884 6959 41893
rect 7285 41833 7341 41842
rect 7681 41898 7737 41907
rect 7681 41833 7737 41842
rect 6903 41819 6959 41828
rect 6046 41526 6102 41535
rect 6046 41461 6102 41470
rect 6471 41526 6527 41535
rect 6471 41461 6527 41470
rect 6903 41526 6959 41535
rect 6903 41461 6959 41470
rect 7285 41503 7341 41512
rect 7285 41438 7341 41447
rect 7681 41503 7737 41512
rect 7681 41438 7737 41447
rect 6046 41152 6102 41161
rect 7285 41108 7341 41117
rect 6046 41087 6102 41096
rect 6471 41094 6527 41103
rect 6471 41029 6527 41038
rect 6903 41094 6959 41103
rect 7285 41043 7341 41052
rect 7681 41108 7737 41117
rect 7681 41043 7737 41052
rect 6903 41029 6959 41038
rect 6046 40736 6102 40745
rect 6046 40671 6102 40680
rect 6471 40736 6527 40745
rect 6471 40671 6527 40680
rect 6903 40736 6959 40745
rect 6903 40671 6959 40680
rect 7285 40713 7341 40722
rect 7285 40648 7341 40657
rect 7681 40713 7737 40722
rect 7681 40648 7737 40657
rect 6046 40362 6102 40371
rect 7285 40318 7341 40327
rect 6046 40297 6102 40306
rect 6471 40304 6527 40313
rect 6471 40239 6527 40248
rect 6903 40304 6959 40313
rect 7285 40253 7341 40262
rect 7681 40318 7737 40327
rect 7681 40253 7737 40262
rect 6903 40239 6959 40248
rect 6046 39946 6102 39955
rect 6046 39881 6102 39890
rect 6471 39946 6527 39955
rect 6471 39881 6527 39890
rect 6903 39946 6959 39955
rect 6903 39881 6959 39890
rect 7285 39923 7341 39932
rect 7285 39858 7341 39867
rect 7681 39923 7737 39932
rect 7681 39858 7737 39867
rect 6046 39572 6102 39581
rect 7285 39528 7341 39537
rect 6046 39507 6102 39516
rect 6471 39514 6527 39523
rect 6471 39449 6527 39458
rect 6903 39514 6959 39523
rect 7285 39463 7341 39472
rect 7681 39528 7737 39537
rect 7681 39463 7737 39472
rect 6903 39449 6959 39458
rect 6046 39156 6102 39165
rect 6046 39091 6102 39100
rect 6471 39156 6527 39165
rect 6471 39091 6527 39100
rect 6903 39156 6959 39165
rect 6903 39091 6959 39100
rect 7285 39133 7341 39142
rect 7285 39068 7341 39077
rect 7681 39133 7737 39142
rect 7681 39068 7737 39077
rect 6046 38782 6102 38791
rect 7285 38738 7341 38747
rect 6046 38717 6102 38726
rect 6471 38724 6527 38733
rect 6471 38659 6527 38668
rect 6903 38724 6959 38733
rect 7285 38673 7341 38682
rect 7681 38738 7737 38747
rect 7681 38673 7737 38682
rect 6903 38659 6959 38668
rect 6046 38366 6102 38375
rect 6046 38301 6102 38310
rect 6471 38366 6527 38375
rect 6471 38301 6527 38310
rect 6903 38366 6959 38375
rect 6903 38301 6959 38310
rect 7285 38343 7341 38352
rect 7285 38278 7341 38287
rect 7681 38343 7737 38352
rect 7681 38278 7737 38287
rect 6046 37992 6102 38001
rect 7285 37948 7341 37957
rect 6046 37927 6102 37936
rect 6471 37934 6527 37943
rect 6471 37869 6527 37878
rect 6903 37934 6959 37943
rect 7285 37883 7341 37892
rect 7681 37948 7737 37957
rect 7681 37883 7737 37892
rect 6903 37869 6959 37878
rect 6046 37576 6102 37585
rect 6046 37511 6102 37520
rect 6471 37576 6527 37585
rect 6471 37511 6527 37520
rect 6903 37576 6959 37585
rect 6903 37511 6959 37520
rect 7285 37553 7341 37562
rect 7285 37488 7341 37497
rect 7681 37553 7737 37562
rect 7681 37488 7737 37497
rect 6046 37202 6102 37211
rect 7285 37158 7341 37167
rect 6046 37137 6102 37146
rect 6471 37144 6527 37153
rect 6471 37079 6527 37088
rect 6903 37144 6959 37153
rect 7285 37093 7341 37102
rect 7681 37158 7737 37167
rect 7681 37093 7737 37102
rect 6903 37079 6959 37088
rect 6046 36786 6102 36795
rect 6046 36721 6102 36730
rect 6471 36786 6527 36795
rect 6471 36721 6527 36730
rect 6903 36786 6959 36795
rect 6903 36721 6959 36730
rect 7285 36763 7341 36772
rect 7285 36698 7341 36707
rect 7681 36763 7737 36772
rect 7681 36698 7737 36707
rect 6046 36412 6102 36421
rect 7285 36368 7341 36377
rect 6046 36347 6102 36356
rect 6471 36354 6527 36363
rect 6471 36289 6527 36298
rect 6903 36354 6959 36363
rect 7285 36303 7341 36312
rect 7681 36368 7737 36377
rect 7681 36303 7737 36312
rect 6903 36289 6959 36298
rect 6046 35996 6102 36005
rect 6046 35931 6102 35940
rect 6471 35996 6527 36005
rect 6471 35931 6527 35940
rect 6903 35996 6959 36005
rect 6903 35931 6959 35940
rect 7285 35973 7341 35982
rect 7285 35908 7341 35917
rect 7681 35973 7737 35982
rect 7681 35908 7737 35917
rect 6046 35622 6102 35631
rect 7285 35578 7341 35587
rect 6046 35557 6102 35566
rect 6471 35564 6527 35573
rect 6471 35499 6527 35508
rect 6903 35564 6959 35573
rect 7285 35513 7341 35522
rect 7681 35578 7737 35587
rect 7681 35513 7737 35522
rect 6903 35499 6959 35508
rect 6046 35206 6102 35215
rect 6046 35141 6102 35150
rect 6471 35206 6527 35215
rect 6471 35141 6527 35150
rect 6903 35206 6959 35215
rect 6903 35141 6959 35150
rect 7285 35183 7341 35192
rect 7285 35118 7341 35127
rect 7681 35183 7737 35192
rect 7681 35118 7737 35127
rect 6046 34832 6102 34841
rect 7285 34788 7341 34797
rect 6046 34767 6102 34776
rect 6471 34774 6527 34783
rect 6471 34709 6527 34718
rect 6903 34774 6959 34783
rect 7285 34723 7341 34732
rect 7681 34788 7737 34797
rect 7681 34723 7737 34732
rect 6903 34709 6959 34718
rect 6046 34416 6102 34425
rect 6046 34351 6102 34360
rect 6471 34416 6527 34425
rect 6471 34351 6527 34360
rect 6903 34416 6959 34425
rect 6903 34351 6959 34360
rect 7285 34393 7341 34402
rect 7285 34328 7341 34337
rect 7681 34393 7737 34402
rect 7681 34328 7737 34337
rect 6046 34042 6102 34051
rect 7285 33998 7341 34007
rect 6046 33977 6102 33986
rect 6471 33984 6527 33993
rect 6471 33919 6527 33928
rect 6903 33984 6959 33993
rect 7285 33933 7341 33942
rect 7681 33998 7737 34007
rect 7681 33933 7737 33942
rect 6903 33919 6959 33928
rect 6046 33626 6102 33635
rect 6046 33561 6102 33570
rect 6471 33626 6527 33635
rect 6471 33561 6527 33570
rect 6903 33626 6959 33635
rect 6903 33561 6959 33570
rect 7285 33603 7341 33612
rect 7285 33538 7341 33547
rect 7681 33603 7737 33612
rect 7681 33538 7737 33547
rect 6046 33252 6102 33261
rect 7285 33208 7341 33217
rect 6046 33187 6102 33196
rect 6471 33194 6527 33203
rect 6471 33129 6527 33138
rect 6903 33194 6959 33203
rect 7285 33143 7341 33152
rect 7681 33208 7737 33217
rect 7681 33143 7737 33152
rect 6903 33129 6959 33138
rect 6046 32836 6102 32845
rect 6046 32771 6102 32780
rect 6471 32836 6527 32845
rect 6471 32771 6527 32780
rect 6903 32836 6959 32845
rect 6903 32771 6959 32780
rect 7285 32813 7341 32822
rect 7285 32748 7341 32757
rect 7681 32813 7737 32822
rect 7681 32748 7737 32757
rect 6046 32462 6102 32471
rect 7285 32418 7341 32427
rect 6046 32397 6102 32406
rect 6471 32404 6527 32413
rect 6471 32339 6527 32348
rect 6903 32404 6959 32413
rect 7285 32353 7341 32362
rect 7681 32418 7737 32427
rect 7681 32353 7737 32362
rect 6903 32339 6959 32348
rect 6046 32046 6102 32055
rect 6046 31981 6102 31990
rect 6471 32046 6527 32055
rect 6471 31981 6527 31990
rect 6903 32046 6959 32055
rect 6903 31981 6959 31990
rect 7285 32023 7341 32032
rect 7285 31958 7341 31967
rect 7681 32023 7737 32032
rect 7681 31958 7737 31967
rect 6046 31672 6102 31681
rect 7285 31628 7341 31637
rect 6046 31607 6102 31616
rect 6471 31614 6527 31623
rect 6471 31549 6527 31558
rect 6903 31614 6959 31623
rect 7285 31563 7341 31572
rect 7681 31628 7737 31637
rect 7681 31563 7737 31572
rect 6903 31549 6959 31558
rect 6046 31256 6102 31265
rect 6046 31191 6102 31200
rect 6471 31256 6527 31265
rect 6471 31191 6527 31200
rect 6903 31256 6959 31265
rect 6903 31191 6959 31200
rect 7285 31233 7341 31242
rect 7285 31168 7341 31177
rect 7681 31233 7737 31242
rect 7681 31168 7737 31177
rect 6046 30882 6102 30891
rect 7285 30838 7341 30847
rect 6046 30817 6102 30826
rect 6471 30824 6527 30833
rect 6471 30759 6527 30768
rect 6903 30824 6959 30833
rect 7285 30773 7341 30782
rect 7681 30838 7737 30847
rect 7681 30773 7737 30782
rect 6903 30759 6959 30768
rect 6046 30466 6102 30475
rect 6046 30401 6102 30410
rect 6471 30466 6527 30475
rect 6471 30401 6527 30410
rect 6903 30466 6959 30475
rect 6903 30401 6959 30410
rect 7285 30443 7341 30452
rect 7285 30378 7341 30387
rect 7681 30443 7737 30452
rect 7681 30378 7737 30387
rect 6046 30092 6102 30101
rect 7285 30048 7341 30057
rect 6046 30027 6102 30036
rect 6471 30034 6527 30043
rect 6471 29969 6527 29978
rect 6903 30034 6959 30043
rect 7285 29983 7341 29992
rect 7681 30048 7737 30057
rect 7681 29983 7737 29992
rect 6903 29969 6959 29978
rect 6046 29676 6102 29685
rect 6046 29611 6102 29620
rect 6471 29676 6527 29685
rect 6471 29611 6527 29620
rect 6903 29676 6959 29685
rect 6903 29611 6959 29620
rect 7285 29653 7341 29662
rect 7285 29588 7341 29597
rect 7681 29653 7737 29662
rect 7681 29588 7737 29597
rect 6046 29302 6102 29311
rect 7285 29258 7341 29267
rect 6046 29237 6102 29246
rect 6471 29244 6527 29253
rect 6471 29179 6527 29188
rect 6903 29244 6959 29253
rect 7285 29193 7341 29202
rect 7681 29258 7737 29267
rect 7681 29193 7737 29202
rect 6903 29179 6959 29188
rect 6046 28886 6102 28895
rect 6046 28821 6102 28830
rect 6471 28886 6527 28895
rect 6471 28821 6527 28830
rect 6903 28886 6959 28895
rect 6903 28821 6959 28830
rect 7285 28863 7341 28872
rect 7285 28798 7341 28807
rect 7681 28863 7737 28872
rect 7681 28798 7737 28807
rect 6046 28512 6102 28521
rect 7285 28468 7341 28477
rect 6046 28447 6102 28456
rect 6471 28454 6527 28463
rect 6471 28389 6527 28398
rect 6903 28454 6959 28463
rect 7285 28403 7341 28412
rect 7681 28468 7737 28477
rect 7681 28403 7737 28412
rect 6903 28389 6959 28398
rect 6046 28096 6102 28105
rect 6046 28031 6102 28040
rect 6471 28096 6527 28105
rect 6471 28031 6527 28040
rect 6903 28096 6959 28105
rect 6903 28031 6959 28040
rect 7285 28073 7341 28082
rect 7285 28008 7341 28017
rect 7681 28073 7737 28082
rect 7681 28008 7737 28017
rect 6046 27722 6102 27731
rect 7285 27678 7341 27687
rect 6046 27657 6102 27666
rect 6471 27664 6527 27673
rect 6471 27599 6527 27608
rect 6903 27664 6959 27673
rect 7285 27613 7341 27622
rect 7681 27678 7737 27687
rect 7681 27613 7737 27622
rect 6903 27599 6959 27608
rect 6046 27306 6102 27315
rect 6046 27241 6102 27250
rect 6471 27306 6527 27315
rect 6471 27241 6527 27250
rect 6903 27306 6959 27315
rect 6903 27241 6959 27250
rect 7285 27283 7341 27292
rect 7285 27218 7341 27227
rect 7681 27283 7737 27292
rect 7681 27218 7737 27227
rect 6046 26932 6102 26941
rect 7285 26888 7341 26897
rect 6046 26867 6102 26876
rect 6471 26874 6527 26883
rect 6471 26809 6527 26818
rect 6903 26874 6959 26883
rect 7285 26823 7341 26832
rect 7681 26888 7737 26897
rect 7681 26823 7737 26832
rect 6903 26809 6959 26818
rect 6046 26516 6102 26525
rect 6046 26451 6102 26460
rect 6471 26516 6527 26525
rect 6471 26451 6527 26460
rect 6903 26516 6959 26525
rect 6903 26451 6959 26460
rect 7285 26493 7341 26502
rect 7285 26428 7341 26437
rect 7681 26493 7737 26502
rect 7681 26428 7737 26437
rect 6046 26142 6102 26151
rect 7285 26098 7341 26107
rect 6046 26077 6102 26086
rect 6471 26084 6527 26093
rect 6471 26019 6527 26028
rect 6903 26084 6959 26093
rect 7285 26033 7341 26042
rect 7681 26098 7737 26107
rect 7681 26033 7737 26042
rect 6903 26019 6959 26028
rect 6046 25726 6102 25735
rect 6046 25661 6102 25670
rect 6471 25726 6527 25735
rect 6471 25661 6527 25670
rect 6903 25726 6959 25735
rect 6903 25661 6959 25670
rect 7285 25703 7341 25712
rect 7285 25638 7341 25647
rect 7681 25703 7737 25712
rect 7681 25638 7737 25647
rect 6046 25352 6102 25361
rect 7285 25308 7341 25317
rect 6046 25287 6102 25296
rect 6471 25294 6527 25303
rect 6471 25229 6527 25238
rect 6903 25294 6959 25303
rect 7285 25243 7341 25252
rect 7681 25308 7737 25317
rect 7681 25243 7737 25252
rect 6903 25229 6959 25238
rect 6046 24936 6102 24945
rect 6046 24871 6102 24880
rect 6471 24936 6527 24945
rect 6471 24871 6527 24880
rect 6903 24936 6959 24945
rect 6903 24871 6959 24880
rect 7285 24913 7341 24922
rect 7285 24848 7341 24857
rect 7681 24913 7737 24922
rect 7681 24848 7737 24857
rect 6046 24562 6102 24571
rect 7285 24518 7341 24527
rect 6046 24497 6102 24506
rect 6471 24504 6527 24513
rect 6471 24439 6527 24448
rect 6903 24504 6959 24513
rect 7285 24453 7341 24462
rect 7681 24518 7737 24527
rect 7681 24453 7737 24462
rect 6903 24439 6959 24448
rect 6046 24146 6102 24155
rect 6046 24081 6102 24090
rect 6471 24146 6527 24155
rect 6471 24081 6527 24090
rect 6903 24146 6959 24155
rect 6903 24081 6959 24090
rect 7285 24123 7341 24132
rect 7285 24058 7341 24067
rect 7681 24123 7737 24132
rect 7681 24058 7737 24067
rect 6046 23772 6102 23781
rect 7285 23728 7341 23737
rect 6046 23707 6102 23716
rect 6471 23714 6527 23723
rect 6471 23649 6527 23658
rect 6903 23714 6959 23723
rect 7285 23663 7341 23672
rect 7681 23728 7737 23737
rect 7681 23663 7737 23672
rect 6903 23649 6959 23658
rect 6046 23356 6102 23365
rect 6046 23291 6102 23300
rect 6471 23356 6527 23365
rect 6471 23291 6527 23300
rect 6903 23356 6959 23365
rect 6903 23291 6959 23300
rect 7285 23333 7341 23342
rect 7285 23268 7341 23277
rect 7681 23333 7737 23342
rect 7681 23268 7737 23277
rect 6046 22982 6102 22991
rect 7285 22938 7341 22947
rect 6046 22917 6102 22926
rect 6471 22924 6527 22933
rect 6471 22859 6527 22868
rect 6903 22924 6959 22933
rect 7285 22873 7341 22882
rect 7681 22938 7737 22947
rect 7681 22873 7737 22882
rect 6903 22859 6959 22868
rect 6046 22566 6102 22575
rect 6046 22501 6102 22510
rect 6471 22566 6527 22575
rect 6471 22501 6527 22510
rect 6903 22566 6959 22575
rect 6903 22501 6959 22510
rect 7285 22543 7341 22552
rect 7285 22478 7341 22487
rect 7681 22543 7737 22552
rect 7681 22478 7737 22487
rect 6046 22192 6102 22201
rect 7285 22148 7341 22157
rect 6046 22127 6102 22136
rect 6471 22134 6527 22143
rect 6471 22069 6527 22078
rect 6903 22134 6959 22143
rect 7285 22083 7341 22092
rect 7681 22148 7737 22157
rect 7681 22083 7737 22092
rect 6903 22069 6959 22078
rect 6046 21776 6102 21785
rect 6046 21711 6102 21720
rect 6471 21776 6527 21785
rect 6471 21711 6527 21720
rect 6903 21776 6959 21785
rect 6903 21711 6959 21720
rect 7285 21753 7341 21762
rect 7285 21688 7341 21697
rect 7681 21753 7737 21762
rect 7681 21688 7737 21697
rect 6046 21402 6102 21411
rect 7285 21358 7341 21367
rect 6046 21337 6102 21346
rect 6471 21344 6527 21353
rect 6471 21279 6527 21288
rect 6903 21344 6959 21353
rect 7285 21293 7341 21302
rect 7681 21358 7737 21367
rect 7681 21293 7737 21302
rect 6903 21279 6959 21288
rect 6046 20986 6102 20995
rect 6046 20921 6102 20930
rect 6471 20986 6527 20995
rect 6471 20921 6527 20930
rect 6903 20986 6959 20995
rect 6903 20921 6959 20930
rect 7285 20963 7341 20972
rect 7285 20898 7341 20907
rect 7681 20963 7737 20972
rect 7681 20898 7737 20907
rect 6046 20612 6102 20621
rect 7285 20568 7341 20577
rect 6046 20547 6102 20556
rect 6471 20554 6527 20563
rect 6471 20489 6527 20498
rect 6903 20554 6959 20563
rect 7285 20503 7341 20512
rect 7681 20568 7737 20577
rect 7681 20503 7737 20512
rect 6903 20489 6959 20498
rect 6046 20196 6102 20205
rect 6046 20131 6102 20140
rect 6471 20196 6527 20205
rect 6471 20131 6527 20140
rect 6903 20196 6959 20205
rect 6903 20131 6959 20140
rect 7285 20173 7341 20182
rect 7285 20108 7341 20117
rect 7681 20173 7737 20182
rect 7681 20108 7737 20117
rect 6046 19822 6102 19831
rect 7285 19778 7341 19787
rect 6046 19757 6102 19766
rect 6471 19764 6527 19773
rect 6471 19699 6527 19708
rect 6903 19764 6959 19773
rect 7285 19713 7341 19722
rect 7681 19778 7737 19787
rect 7681 19713 7737 19722
rect 6903 19699 6959 19708
rect 6046 19406 6102 19415
rect 6046 19341 6102 19350
rect 6471 19406 6527 19415
rect 6471 19341 6527 19350
rect 6903 19406 6959 19415
rect 6903 19341 6959 19350
rect 7285 19383 7341 19392
rect 7285 19318 7341 19327
rect 7681 19383 7737 19392
rect 7681 19318 7737 19327
rect 6046 19032 6102 19041
rect 7285 18988 7341 18997
rect 6046 18967 6102 18976
rect 6471 18974 6527 18983
rect 6471 18909 6527 18918
rect 6903 18974 6959 18983
rect 7285 18923 7341 18932
rect 7681 18988 7737 18997
rect 7681 18923 7737 18932
rect 6903 18909 6959 18918
rect 6046 18616 6102 18625
rect 6046 18551 6102 18560
rect 6471 18616 6527 18625
rect 6471 18551 6527 18560
rect 6903 18616 6959 18625
rect 6903 18551 6959 18560
rect 7285 18593 7341 18602
rect 7285 18528 7341 18537
rect 7681 18593 7737 18602
rect 7681 18528 7737 18537
rect 6046 18242 6102 18251
rect 7285 18198 7341 18207
rect 6046 18177 6102 18186
rect 6471 18184 6527 18193
rect 6471 18119 6527 18128
rect 6903 18184 6959 18193
rect 7285 18133 7341 18142
rect 7681 18198 7737 18207
rect 7681 18133 7737 18142
rect 6903 18119 6959 18128
rect 6046 17826 6102 17835
rect 6046 17761 6102 17770
rect 6471 17826 6527 17835
rect 6471 17761 6527 17770
rect 6903 17826 6959 17835
rect 6903 17761 6959 17770
rect 7285 17803 7341 17812
rect 7285 17738 7341 17747
rect 7681 17803 7737 17812
rect 7681 17738 7737 17747
rect 6046 17452 6102 17461
rect 7285 17408 7341 17417
rect 6046 17387 6102 17396
rect 6471 17394 6527 17403
rect 6471 17329 6527 17338
rect 6903 17394 6959 17403
rect 7285 17343 7341 17352
rect 7681 17408 7737 17417
rect 7681 17343 7737 17352
rect 6903 17329 6959 17338
rect 6046 17036 6102 17045
rect 6046 16971 6102 16980
rect 6471 17036 6527 17045
rect 6471 16971 6527 16980
rect 6903 17036 6959 17045
rect 6903 16971 6959 16980
rect 7285 17013 7341 17022
rect 7285 16948 7341 16957
rect 7681 17013 7737 17022
rect 7681 16948 7737 16957
rect 6046 16662 6102 16671
rect 7285 16618 7341 16627
rect 6046 16597 6102 16606
rect 6471 16604 6527 16613
rect 6471 16539 6527 16548
rect 6903 16604 6959 16613
rect 7285 16553 7341 16562
rect 7681 16618 7737 16627
rect 7681 16553 7737 16562
rect 6903 16539 6959 16548
rect 6046 16246 6102 16255
rect 6046 16181 6102 16190
rect 6471 16246 6527 16255
rect 6471 16181 6527 16190
rect 6903 16246 6959 16255
rect 6903 16181 6959 16190
rect 7285 16223 7341 16232
rect 7285 16158 7341 16167
rect 7681 16223 7737 16232
rect 7681 16158 7737 16167
rect 6046 15872 6102 15881
rect 7285 15828 7341 15837
rect 6046 15807 6102 15816
rect 6471 15814 6527 15823
rect 6471 15749 6527 15758
rect 6903 15814 6959 15823
rect 7285 15763 7341 15772
rect 7681 15828 7737 15837
rect 7681 15763 7737 15772
rect 6903 15749 6959 15758
rect 6046 15456 6102 15465
rect 6046 15391 6102 15400
rect 6471 15456 6527 15465
rect 6471 15391 6527 15400
rect 6903 15456 6959 15465
rect 6903 15391 6959 15400
rect 7285 15433 7341 15442
rect 7285 15368 7341 15377
rect 7681 15433 7737 15442
rect 7681 15368 7737 15377
rect 6046 15082 6102 15091
rect 7285 15038 7341 15047
rect 6046 15017 6102 15026
rect 6471 15024 6527 15033
rect 6471 14959 6527 14968
rect 6903 15024 6959 15033
rect 7285 14973 7341 14982
rect 7681 15038 7737 15047
rect 7681 14973 7737 14982
rect 6903 14959 6959 14968
rect 6046 14666 6102 14675
rect 6046 14601 6102 14610
rect 6471 14666 6527 14675
rect 6471 14601 6527 14610
rect 6903 14666 6959 14675
rect 6903 14601 6959 14610
rect 7285 14643 7341 14652
rect 7285 14578 7341 14587
rect 7681 14643 7737 14652
rect 7681 14578 7737 14587
rect 6046 14292 6102 14301
rect 7285 14248 7341 14257
rect 6046 14227 6102 14236
rect 6471 14234 6527 14243
rect 6471 14169 6527 14178
rect 6903 14234 6959 14243
rect 7285 14183 7341 14192
rect 7681 14248 7737 14257
rect 7681 14183 7737 14192
rect 6903 14169 6959 14178
rect 6046 13876 6102 13885
rect 6046 13811 6102 13820
rect 6471 13876 6527 13885
rect 6471 13811 6527 13820
rect 6903 13876 6959 13885
rect 6903 13811 6959 13820
rect 7285 13853 7341 13862
rect 7285 13788 7341 13797
rect 7681 13853 7737 13862
rect 7681 13788 7737 13797
rect 6046 13502 6102 13511
rect 7285 13458 7341 13467
rect 6046 13437 6102 13446
rect 6471 13444 6527 13453
rect 6471 13379 6527 13388
rect 6903 13444 6959 13453
rect 7285 13393 7341 13402
rect 7681 13458 7737 13467
rect 7681 13393 7737 13402
rect 6903 13379 6959 13388
rect 6046 13086 6102 13095
rect 6046 13021 6102 13030
rect 6471 13086 6527 13095
rect 6471 13021 6527 13030
rect 6903 13086 6959 13095
rect 6903 13021 6959 13030
rect 7285 13063 7341 13072
rect 7285 12998 7341 13007
rect 7681 13063 7737 13072
rect 7681 12998 7737 13007
rect 6046 12712 6102 12721
rect 7285 12668 7341 12677
rect 6046 12647 6102 12656
rect 6471 12654 6527 12663
rect 6471 12589 6527 12598
rect 6903 12654 6959 12663
rect 7285 12603 7341 12612
rect 7681 12668 7737 12677
rect 7681 12603 7737 12612
rect 6903 12589 6959 12598
rect 6046 12296 6102 12305
rect 6046 12231 6102 12240
rect 6471 12296 6527 12305
rect 6471 12231 6527 12240
rect 6903 12296 6959 12305
rect 6903 12231 6959 12240
rect 7285 12273 7341 12282
rect 7285 12208 7341 12217
rect 7681 12273 7737 12282
rect 7681 12208 7737 12217
rect 6046 11922 6102 11931
rect 7285 11878 7341 11887
rect 6046 11857 6102 11866
rect 6471 11864 6527 11873
rect 6471 11799 6527 11808
rect 6903 11864 6959 11873
rect 7285 11813 7341 11822
rect 7681 11878 7737 11887
rect 7681 11813 7737 11822
rect 6903 11799 6959 11808
rect 6046 11506 6102 11515
rect 6046 11441 6102 11450
rect 6471 11506 6527 11515
rect 6471 11441 6527 11450
rect 6903 11506 6959 11515
rect 6903 11441 6959 11450
rect 7285 11483 7341 11492
rect 7285 11418 7341 11427
rect 7681 11483 7737 11492
rect 7681 11418 7737 11427
rect 6046 11132 6102 11141
rect 7285 11088 7341 11097
rect 6046 11067 6102 11076
rect 6471 11074 6527 11083
rect 6471 11009 6527 11018
rect 6903 11074 6959 11083
rect 7285 11023 7341 11032
rect 7681 11088 7737 11097
rect 7681 11023 7737 11032
rect 6903 11009 6959 11018
rect 6046 10716 6102 10725
rect 6046 10651 6102 10660
rect 6471 10716 6527 10725
rect 6471 10651 6527 10660
rect 6903 10716 6959 10725
rect 6903 10651 6959 10660
rect 7285 10693 7341 10702
rect 7285 10628 7341 10637
rect 7681 10693 7737 10702
rect 7681 10628 7737 10637
rect 6046 10342 6102 10351
rect 7285 10298 7341 10307
rect 6046 10277 6102 10286
rect 6471 10284 6527 10293
rect 6471 10219 6527 10228
rect 6903 10284 6959 10293
rect 7285 10233 7341 10242
rect 7681 10298 7737 10307
rect 7681 10233 7737 10242
rect 6903 10219 6959 10228
rect 6046 9926 6102 9935
rect 6046 9861 6102 9870
rect 6471 9926 6527 9935
rect 6471 9861 6527 9870
rect 6903 9926 6959 9935
rect 6903 9861 6959 9870
rect 7285 9903 7341 9912
rect 7285 9838 7341 9847
rect 7681 9903 7737 9912
rect 7681 9838 7737 9847
rect 6046 9552 6102 9561
rect 7285 9508 7341 9517
rect 6046 9487 6102 9496
rect 6471 9494 6527 9503
rect 6471 9429 6527 9438
rect 6903 9494 6959 9503
rect 7285 9443 7341 9452
rect 7681 9508 7737 9517
rect 7681 9443 7737 9452
rect 6903 9429 6959 9438
rect 6046 9136 6102 9145
rect 6046 9071 6102 9080
rect 6471 9136 6527 9145
rect 6471 9071 6527 9080
rect 6903 9136 6959 9145
rect 6903 9071 6959 9080
rect 7285 9113 7341 9122
rect 7285 9048 7341 9057
rect 7681 9113 7737 9122
rect 7681 9048 7737 9057
rect 6046 8762 6102 8771
rect 7285 8718 7341 8727
rect 6046 8697 6102 8706
rect 6471 8704 6527 8713
rect 6471 8639 6527 8648
rect 6903 8704 6959 8713
rect 7285 8653 7341 8662
rect 7681 8718 7737 8727
rect 7681 8653 7737 8662
rect 6903 8639 6959 8648
rect 6046 8346 6102 8355
rect 6046 8281 6102 8290
rect 6471 8346 6527 8355
rect 6471 8281 6527 8290
rect 6903 8346 6959 8355
rect 6903 8281 6959 8290
rect 7285 8323 7341 8332
rect 7285 8258 7341 8267
rect 7681 8323 7737 8332
rect 7681 8258 7737 8267
rect 6046 7972 6102 7981
rect 7285 7928 7341 7937
rect 6046 7907 6102 7916
rect 6471 7914 6527 7923
rect 6471 7849 6527 7858
rect 6903 7914 6959 7923
rect 7285 7863 7341 7872
rect 7681 7928 7737 7937
rect 7681 7863 7737 7872
rect 6903 7849 6959 7858
rect 4417 7806 4469 7812
rect 4469 7766 4541 7794
rect 4417 7748 4469 7754
rect 4513 7519 4541 7766
rect 6046 7556 6102 7565
rect 5705 7519 5711 7531
rect 4513 7491 5711 7519
rect 5705 7479 5711 7491
rect 5763 7479 5769 7531
rect 6046 7491 6102 7500
rect 6471 7556 6527 7565
rect 6471 7491 6527 7500
rect 6903 7556 6959 7565
rect 6903 7491 6959 7500
rect 7285 7533 7341 7542
rect 7285 7468 7341 7477
rect 7681 7533 7737 7542
rect 7681 7468 7737 7477
rect 4417 7256 4469 7262
rect 4469 7216 4541 7244
rect 4417 7198 4469 7204
rect 4513 7124 4541 7216
rect 6046 7182 6102 7191
rect 5625 7124 5631 7136
rect 4513 7096 5631 7124
rect 5625 7084 5631 7096
rect 5683 7084 5689 7136
rect 7285 7138 7341 7147
rect 6046 7117 6102 7126
rect 6471 7124 6527 7133
rect 6471 7059 6527 7068
rect 6903 7124 6959 7133
rect 7285 7073 7341 7082
rect 7681 7138 7737 7147
rect 7681 7073 7737 7082
rect 6903 7059 6959 7068
rect 4417 7016 4469 7022
rect 4469 6976 4541 7004
rect 4417 6958 4469 6964
rect 4513 6729 4541 6976
rect 6046 6766 6102 6775
rect 5545 6729 5551 6741
rect 4513 6701 5551 6729
rect 5545 6689 5551 6701
rect 5603 6689 5609 6741
rect 6046 6701 6102 6710
rect 6471 6766 6527 6775
rect 6471 6701 6527 6710
rect 6903 6766 6959 6775
rect 6903 6701 6959 6710
rect 7285 6743 7341 6752
rect 7285 6678 7341 6687
rect 7681 6743 7737 6752
rect 7681 6678 7737 6687
rect 4417 6466 4469 6472
rect 4469 6426 4541 6454
rect 4417 6408 4469 6414
rect 4513 6334 4541 6426
rect 6046 6392 6102 6401
rect 5465 6334 5471 6346
rect 4513 6306 5471 6334
rect 5465 6294 5471 6306
rect 5523 6294 5529 6346
rect 7285 6348 7341 6357
rect 6046 6327 6102 6336
rect 6471 6334 6527 6343
rect 6471 6269 6527 6278
rect 6903 6334 6959 6343
rect 7285 6283 7341 6292
rect 7681 6348 7737 6357
rect 7681 6283 7737 6292
rect 6903 6269 6959 6278
rect 4417 6226 4469 6232
rect 4469 6186 4541 6214
rect 4417 6168 4469 6174
rect 4513 5939 4541 6186
rect 6046 5976 6102 5985
rect 5385 5939 5391 5951
rect 4513 5911 5391 5939
rect 5385 5899 5391 5911
rect 5443 5899 5449 5951
rect 6046 5911 6102 5920
rect 6471 5976 6527 5985
rect 6471 5911 6527 5920
rect 6903 5976 6959 5985
rect 6903 5911 6959 5920
rect 7285 5953 7341 5962
rect 7285 5888 7341 5897
rect 7681 5953 7737 5962
rect 7681 5888 7737 5897
rect 4417 5676 4469 5682
rect 4469 5636 4541 5664
rect 4417 5618 4469 5624
rect 4513 5544 4541 5636
rect 6046 5602 6102 5611
rect 5305 5544 5311 5556
rect 4513 5516 5311 5544
rect 5305 5504 5311 5516
rect 5363 5504 5369 5556
rect 7285 5558 7341 5567
rect 6046 5537 6102 5546
rect 6471 5544 6527 5553
rect 6471 5479 6527 5488
rect 6903 5544 6959 5553
rect 7285 5493 7341 5502
rect 7681 5558 7737 5567
rect 7681 5493 7737 5502
rect 6903 5479 6959 5488
rect 4417 5436 4469 5442
rect 4469 5396 4541 5424
rect 4417 5378 4469 5384
rect 4513 5149 4541 5396
rect 6046 5186 6102 5195
rect 5225 5149 5231 5161
rect 4513 5121 5231 5149
rect 5225 5109 5231 5121
rect 5283 5109 5289 5161
rect 6046 5121 6102 5130
rect 6471 5186 6527 5195
rect 6471 5121 6527 5130
rect 6903 5186 6959 5195
rect 6903 5121 6959 5130
rect 7285 5163 7341 5172
rect 7285 5098 7341 5107
rect 7681 5163 7737 5172
rect 7681 5098 7737 5107
rect 4417 4886 4469 4892
rect 4469 4846 4541 4874
rect 4417 4828 4469 4834
rect 4513 4754 4541 4846
rect 6046 4812 6102 4821
rect 5145 4754 5151 4766
rect 4513 4726 5151 4754
rect 5145 4714 5151 4726
rect 5203 4714 5209 4766
rect 7285 4768 7341 4777
rect 6046 4747 6102 4756
rect 6471 4754 6527 4763
rect 6471 4689 6527 4698
rect 6903 4754 6959 4763
rect 7285 4703 7341 4712
rect 7681 4768 7737 4777
rect 7681 4703 7737 4712
rect 6903 4689 6959 4698
rect 6046 4396 6102 4405
rect 6046 4331 6102 4340
rect 6471 4396 6527 4405
rect 6471 4331 6527 4340
rect 6903 4396 6959 4405
rect 6903 4331 6959 4340
rect 7285 4373 7341 4382
rect 7285 4308 7341 4317
rect 7681 4373 7737 4382
rect 7681 4308 7737 4317
rect 6046 4022 6102 4031
rect 7285 3978 7341 3987
rect 6046 3957 6102 3966
rect 6471 3964 6527 3973
rect 6471 3899 6527 3908
rect 6903 3964 6959 3973
rect 7285 3913 7341 3922
rect 7681 3978 7737 3987
rect 7681 3913 7737 3922
rect 6903 3899 6959 3908
rect 4417 3856 4469 3862
rect 4469 3816 4541 3844
rect 4417 3798 4469 3804
rect 4513 3569 4541 3816
rect 6046 3606 6102 3615
rect 5065 3569 5071 3581
rect 4513 3541 5071 3569
rect 5065 3529 5071 3541
rect 5123 3529 5129 3581
rect 6046 3541 6102 3550
rect 6471 3606 6527 3615
rect 6471 3541 6527 3550
rect 6903 3606 6959 3615
rect 6903 3541 6959 3550
rect 7285 3583 7341 3592
rect 7285 3518 7341 3527
rect 7681 3583 7737 3592
rect 7681 3518 7737 3527
rect 4417 3306 4469 3312
rect 4469 3266 4541 3294
rect 4417 3248 4469 3254
rect 4513 3174 4541 3266
rect 6046 3232 6102 3241
rect 4985 3174 4991 3186
rect 4513 3146 4991 3174
rect 4985 3134 4991 3146
rect 5043 3134 5049 3186
rect 7285 3188 7341 3197
rect 6046 3167 6102 3176
rect 6471 3174 6527 3183
rect 6471 3109 6527 3118
rect 6903 3174 6959 3183
rect 7285 3123 7341 3132
rect 7681 3188 7737 3197
rect 7681 3123 7737 3132
rect 6903 3109 6959 3118
rect 4417 3066 4469 3072
rect 4469 3026 4541 3054
rect 4417 3008 4469 3014
rect 4513 2779 4541 3026
rect 6046 2816 6102 2825
rect 4905 2779 4911 2791
rect 4513 2751 4911 2779
rect 4905 2739 4911 2751
rect 4963 2739 4969 2791
rect 6046 2751 6102 2760
rect 6471 2816 6527 2825
rect 6471 2751 6527 2760
rect 6903 2816 6959 2825
rect 6903 2751 6959 2760
rect 7285 2793 7341 2802
rect 7285 2728 7341 2737
rect 7681 2793 7737 2802
rect 7681 2728 7737 2737
rect 4417 2516 4469 2522
rect 4469 2476 4541 2504
rect 4417 2458 4469 2464
rect 4513 2384 4541 2476
rect 6046 2442 6102 2451
rect 4825 2384 4831 2396
rect 4513 2356 4831 2384
rect 4825 2344 4831 2356
rect 4883 2344 4889 2396
rect 7285 2398 7341 2407
rect 6046 2377 6102 2386
rect 6471 2384 6527 2393
rect 6471 2319 6527 2328
rect 6903 2384 6959 2393
rect 7285 2333 7341 2342
rect 7681 2398 7737 2407
rect 7681 2333 7737 2342
rect 6903 2319 6959 2328
rect 6046 2026 6102 2035
rect 6046 1961 6102 1970
rect 6471 2026 6527 2035
rect 6471 1961 6527 1970
rect 6903 2026 6959 2035
rect 6903 1961 6959 1970
rect 7285 2003 7341 2012
rect 7285 1938 7341 1947
rect 7681 2003 7737 2012
rect 7681 1938 7737 1947
rect 6046 1652 6102 1661
rect 7285 1608 7341 1617
rect 6046 1587 6102 1596
rect 6471 1594 6527 1603
rect 6471 1529 6527 1538
rect 6903 1594 6959 1603
rect 7285 1543 7341 1552
rect 7681 1608 7737 1617
rect 7681 1543 7737 1552
rect 6903 1529 6959 1538
rect 4417 1486 4469 1492
rect 4469 1446 4541 1474
rect 4417 1428 4469 1434
rect 4513 1199 4541 1446
rect 6046 1236 6102 1245
rect 4745 1199 4751 1211
rect 4513 1171 4751 1199
rect 4745 1159 4751 1171
rect 4803 1159 4809 1211
rect 6046 1171 6102 1180
rect 6471 1236 6527 1245
rect 6471 1171 6527 1180
rect 6903 1236 6959 1245
rect 6903 1171 6959 1180
rect 7285 1213 7341 1222
rect 7285 1148 7341 1157
rect 7681 1213 7737 1222
rect 7681 1148 7737 1157
rect 4417 936 4469 942
rect 4469 896 4541 924
rect 4417 878 4469 884
rect 4513 804 4541 896
rect 6046 862 6102 871
rect 4665 804 4671 816
rect 4513 776 4671 804
rect 4665 764 4671 776
rect 4723 764 4729 816
rect 7285 818 7341 827
rect 6046 797 6102 806
rect 6471 804 6527 813
rect 6471 739 6527 748
rect 6903 804 6959 813
rect 7285 753 7341 762
rect 7681 818 7737 827
rect 7681 753 7737 762
rect 6903 739 6959 748
rect 4417 696 4469 702
rect 4469 656 4541 684
rect 4417 638 4469 644
rect 4513 409 4541 656
rect 6046 446 6102 455
rect 4585 409 4591 421
rect 4513 381 4591 409
rect 4585 369 4591 381
rect 4643 369 4649 421
rect 6046 381 6102 390
rect 6471 446 6527 455
rect 6471 381 6527 390
rect 6903 446 6959 455
rect 6903 381 6959 390
rect 7285 423 7341 432
rect 7285 358 7341 367
rect 7681 423 7737 432
rect 7681 358 7737 367
rect 4417 146 4469 152
rect 4469 106 4541 134
rect 4417 88 4469 94
rect 4513 26 4541 106
rect 4505 -26 4511 26
rect 4563 -26 4569 26
<< via2 >>
rect 6046 50214 6102 50216
rect 6046 50162 6048 50214
rect 6048 50162 6100 50214
rect 6100 50162 6102 50214
rect 6046 50160 6102 50162
rect 6471 50214 6527 50216
rect 6471 50162 6473 50214
rect 6473 50162 6525 50214
rect 6525 50162 6527 50214
rect 6471 50160 6527 50162
rect 6903 50214 6959 50216
rect 6903 50162 6905 50214
rect 6905 50162 6957 50214
rect 6957 50162 6959 50214
rect 6903 50160 6959 50162
rect 7285 50191 7341 50193
rect 7285 50139 7287 50191
rect 7287 50139 7339 50191
rect 7339 50139 7341 50191
rect 7285 50137 7341 50139
rect 7681 50191 7737 50193
rect 7681 50139 7683 50191
rect 7683 50139 7735 50191
rect 7735 50139 7737 50191
rect 7681 50137 7737 50139
rect 6046 49840 6102 49842
rect 6046 49788 6048 49840
rect 6048 49788 6100 49840
rect 6100 49788 6102 49840
rect 7285 49796 7341 49798
rect 6046 49786 6102 49788
rect 6471 49782 6527 49784
rect 6471 49730 6473 49782
rect 6473 49730 6525 49782
rect 6525 49730 6527 49782
rect 6471 49728 6527 49730
rect 6903 49782 6959 49784
rect 6903 49730 6905 49782
rect 6905 49730 6957 49782
rect 6957 49730 6959 49782
rect 7285 49744 7287 49796
rect 7287 49744 7339 49796
rect 7339 49744 7341 49796
rect 7285 49742 7341 49744
rect 7681 49796 7737 49798
rect 7681 49744 7683 49796
rect 7683 49744 7735 49796
rect 7735 49744 7737 49796
rect 7681 49742 7737 49744
rect 6903 49728 6959 49730
rect 6046 49424 6102 49426
rect 6046 49372 6048 49424
rect 6048 49372 6100 49424
rect 6100 49372 6102 49424
rect 6046 49370 6102 49372
rect 6471 49424 6527 49426
rect 6471 49372 6473 49424
rect 6473 49372 6525 49424
rect 6525 49372 6527 49424
rect 6471 49370 6527 49372
rect 6903 49424 6959 49426
rect 6903 49372 6905 49424
rect 6905 49372 6957 49424
rect 6957 49372 6959 49424
rect 6903 49370 6959 49372
rect 7285 49401 7341 49403
rect 7285 49349 7287 49401
rect 7287 49349 7339 49401
rect 7339 49349 7341 49401
rect 7285 49347 7341 49349
rect 7681 49401 7737 49403
rect 7681 49349 7683 49401
rect 7683 49349 7735 49401
rect 7735 49349 7737 49401
rect 7681 49347 7737 49349
rect 6046 49050 6102 49052
rect 6046 48998 6048 49050
rect 6048 48998 6100 49050
rect 6100 48998 6102 49050
rect 7285 49006 7341 49008
rect 6046 48996 6102 48998
rect 6471 48992 6527 48994
rect 6471 48940 6473 48992
rect 6473 48940 6525 48992
rect 6525 48940 6527 48992
rect 6471 48938 6527 48940
rect 6903 48992 6959 48994
rect 6903 48940 6905 48992
rect 6905 48940 6957 48992
rect 6957 48940 6959 48992
rect 7285 48954 7287 49006
rect 7287 48954 7339 49006
rect 7339 48954 7341 49006
rect 7285 48952 7341 48954
rect 7681 49006 7737 49008
rect 7681 48954 7683 49006
rect 7683 48954 7735 49006
rect 7735 48954 7737 49006
rect 7681 48952 7737 48954
rect 6903 48938 6959 48940
rect 6046 48634 6102 48636
rect 6046 48582 6048 48634
rect 6048 48582 6100 48634
rect 6100 48582 6102 48634
rect 6046 48580 6102 48582
rect 6471 48634 6527 48636
rect 6471 48582 6473 48634
rect 6473 48582 6525 48634
rect 6525 48582 6527 48634
rect 6471 48580 6527 48582
rect 6903 48634 6959 48636
rect 6903 48582 6905 48634
rect 6905 48582 6957 48634
rect 6957 48582 6959 48634
rect 6903 48580 6959 48582
rect 7285 48611 7341 48613
rect 7285 48559 7287 48611
rect 7287 48559 7339 48611
rect 7339 48559 7341 48611
rect 7285 48557 7341 48559
rect 7681 48611 7737 48613
rect 7681 48559 7683 48611
rect 7683 48559 7735 48611
rect 7735 48559 7737 48611
rect 7681 48557 7737 48559
rect 6046 48260 6102 48262
rect 6046 48208 6048 48260
rect 6048 48208 6100 48260
rect 6100 48208 6102 48260
rect 7285 48216 7341 48218
rect 6046 48206 6102 48208
rect 6471 48202 6527 48204
rect 6471 48150 6473 48202
rect 6473 48150 6525 48202
rect 6525 48150 6527 48202
rect 6471 48148 6527 48150
rect 6903 48202 6959 48204
rect 6903 48150 6905 48202
rect 6905 48150 6957 48202
rect 6957 48150 6959 48202
rect 7285 48164 7287 48216
rect 7287 48164 7339 48216
rect 7339 48164 7341 48216
rect 7285 48162 7341 48164
rect 7681 48216 7737 48218
rect 7681 48164 7683 48216
rect 7683 48164 7735 48216
rect 7735 48164 7737 48216
rect 7681 48162 7737 48164
rect 6903 48148 6959 48150
rect 6046 47844 6102 47846
rect 6046 47792 6048 47844
rect 6048 47792 6100 47844
rect 6100 47792 6102 47844
rect 6046 47790 6102 47792
rect 6471 47844 6527 47846
rect 6471 47792 6473 47844
rect 6473 47792 6525 47844
rect 6525 47792 6527 47844
rect 6471 47790 6527 47792
rect 6903 47844 6959 47846
rect 6903 47792 6905 47844
rect 6905 47792 6957 47844
rect 6957 47792 6959 47844
rect 6903 47790 6959 47792
rect 7285 47821 7341 47823
rect 7285 47769 7287 47821
rect 7287 47769 7339 47821
rect 7339 47769 7341 47821
rect 7285 47767 7341 47769
rect 7681 47821 7737 47823
rect 7681 47769 7683 47821
rect 7683 47769 7735 47821
rect 7735 47769 7737 47821
rect 7681 47767 7737 47769
rect 6046 47470 6102 47472
rect 6046 47418 6048 47470
rect 6048 47418 6100 47470
rect 6100 47418 6102 47470
rect 7285 47426 7341 47428
rect 6046 47416 6102 47418
rect 6471 47412 6527 47414
rect 6471 47360 6473 47412
rect 6473 47360 6525 47412
rect 6525 47360 6527 47412
rect 6471 47358 6527 47360
rect 6903 47412 6959 47414
rect 6903 47360 6905 47412
rect 6905 47360 6957 47412
rect 6957 47360 6959 47412
rect 7285 47374 7287 47426
rect 7287 47374 7339 47426
rect 7339 47374 7341 47426
rect 7285 47372 7341 47374
rect 7681 47426 7737 47428
rect 7681 47374 7683 47426
rect 7683 47374 7735 47426
rect 7735 47374 7737 47426
rect 7681 47372 7737 47374
rect 6903 47358 6959 47360
rect 6046 47054 6102 47056
rect 6046 47002 6048 47054
rect 6048 47002 6100 47054
rect 6100 47002 6102 47054
rect 6046 47000 6102 47002
rect 6471 47054 6527 47056
rect 6471 47002 6473 47054
rect 6473 47002 6525 47054
rect 6525 47002 6527 47054
rect 6471 47000 6527 47002
rect 6903 47054 6959 47056
rect 6903 47002 6905 47054
rect 6905 47002 6957 47054
rect 6957 47002 6959 47054
rect 6903 47000 6959 47002
rect 7285 47031 7341 47033
rect 7285 46979 7287 47031
rect 7287 46979 7339 47031
rect 7339 46979 7341 47031
rect 7285 46977 7341 46979
rect 7681 47031 7737 47033
rect 7681 46979 7683 47031
rect 7683 46979 7735 47031
rect 7735 46979 7737 47031
rect 7681 46977 7737 46979
rect 6046 46680 6102 46682
rect 6046 46628 6048 46680
rect 6048 46628 6100 46680
rect 6100 46628 6102 46680
rect 7285 46636 7341 46638
rect 6046 46626 6102 46628
rect 6471 46622 6527 46624
rect 6471 46570 6473 46622
rect 6473 46570 6525 46622
rect 6525 46570 6527 46622
rect 6471 46568 6527 46570
rect 6903 46622 6959 46624
rect 6903 46570 6905 46622
rect 6905 46570 6957 46622
rect 6957 46570 6959 46622
rect 7285 46584 7287 46636
rect 7287 46584 7339 46636
rect 7339 46584 7341 46636
rect 7285 46582 7341 46584
rect 7681 46636 7737 46638
rect 7681 46584 7683 46636
rect 7683 46584 7735 46636
rect 7735 46584 7737 46636
rect 7681 46582 7737 46584
rect 6903 46568 6959 46570
rect 6046 46264 6102 46266
rect 6046 46212 6048 46264
rect 6048 46212 6100 46264
rect 6100 46212 6102 46264
rect 6046 46210 6102 46212
rect 6471 46264 6527 46266
rect 6471 46212 6473 46264
rect 6473 46212 6525 46264
rect 6525 46212 6527 46264
rect 6471 46210 6527 46212
rect 6903 46264 6959 46266
rect 6903 46212 6905 46264
rect 6905 46212 6957 46264
rect 6957 46212 6959 46264
rect 6903 46210 6959 46212
rect 7285 46241 7341 46243
rect 7285 46189 7287 46241
rect 7287 46189 7339 46241
rect 7339 46189 7341 46241
rect 7285 46187 7341 46189
rect 7681 46241 7737 46243
rect 7681 46189 7683 46241
rect 7683 46189 7735 46241
rect 7735 46189 7737 46241
rect 7681 46187 7737 46189
rect 6046 45890 6102 45892
rect 6046 45838 6048 45890
rect 6048 45838 6100 45890
rect 6100 45838 6102 45890
rect 7285 45846 7341 45848
rect 6046 45836 6102 45838
rect 6471 45832 6527 45834
rect 6471 45780 6473 45832
rect 6473 45780 6525 45832
rect 6525 45780 6527 45832
rect 6471 45778 6527 45780
rect 6903 45832 6959 45834
rect 6903 45780 6905 45832
rect 6905 45780 6957 45832
rect 6957 45780 6959 45832
rect 7285 45794 7287 45846
rect 7287 45794 7339 45846
rect 7339 45794 7341 45846
rect 7285 45792 7341 45794
rect 7681 45846 7737 45848
rect 7681 45794 7683 45846
rect 7683 45794 7735 45846
rect 7735 45794 7737 45846
rect 7681 45792 7737 45794
rect 6903 45778 6959 45780
rect 6046 45474 6102 45476
rect 6046 45422 6048 45474
rect 6048 45422 6100 45474
rect 6100 45422 6102 45474
rect 6046 45420 6102 45422
rect 6471 45474 6527 45476
rect 6471 45422 6473 45474
rect 6473 45422 6525 45474
rect 6525 45422 6527 45474
rect 6471 45420 6527 45422
rect 6903 45474 6959 45476
rect 6903 45422 6905 45474
rect 6905 45422 6957 45474
rect 6957 45422 6959 45474
rect 6903 45420 6959 45422
rect 7285 45451 7341 45453
rect 7285 45399 7287 45451
rect 7287 45399 7339 45451
rect 7339 45399 7341 45451
rect 7285 45397 7341 45399
rect 7681 45451 7737 45453
rect 7681 45399 7683 45451
rect 7683 45399 7735 45451
rect 7735 45399 7737 45451
rect 7681 45397 7737 45399
rect 6046 45100 6102 45102
rect 6046 45048 6048 45100
rect 6048 45048 6100 45100
rect 6100 45048 6102 45100
rect 7285 45056 7341 45058
rect 6046 45046 6102 45048
rect 6471 45042 6527 45044
rect 6471 44990 6473 45042
rect 6473 44990 6525 45042
rect 6525 44990 6527 45042
rect 6471 44988 6527 44990
rect 6903 45042 6959 45044
rect 6903 44990 6905 45042
rect 6905 44990 6957 45042
rect 6957 44990 6959 45042
rect 7285 45004 7287 45056
rect 7287 45004 7339 45056
rect 7339 45004 7341 45056
rect 7285 45002 7341 45004
rect 7681 45056 7737 45058
rect 7681 45004 7683 45056
rect 7683 45004 7735 45056
rect 7735 45004 7737 45056
rect 7681 45002 7737 45004
rect 6903 44988 6959 44990
rect 6046 44684 6102 44686
rect 6046 44632 6048 44684
rect 6048 44632 6100 44684
rect 6100 44632 6102 44684
rect 6046 44630 6102 44632
rect 6471 44684 6527 44686
rect 6471 44632 6473 44684
rect 6473 44632 6525 44684
rect 6525 44632 6527 44684
rect 6471 44630 6527 44632
rect 6903 44684 6959 44686
rect 6903 44632 6905 44684
rect 6905 44632 6957 44684
rect 6957 44632 6959 44684
rect 6903 44630 6959 44632
rect 7285 44661 7341 44663
rect 7285 44609 7287 44661
rect 7287 44609 7339 44661
rect 7339 44609 7341 44661
rect 7285 44607 7341 44609
rect 7681 44661 7737 44663
rect 7681 44609 7683 44661
rect 7683 44609 7735 44661
rect 7735 44609 7737 44661
rect 7681 44607 7737 44609
rect 6046 44310 6102 44312
rect 6046 44258 6048 44310
rect 6048 44258 6100 44310
rect 6100 44258 6102 44310
rect 7285 44266 7341 44268
rect 6046 44256 6102 44258
rect 6471 44252 6527 44254
rect 6471 44200 6473 44252
rect 6473 44200 6525 44252
rect 6525 44200 6527 44252
rect 6471 44198 6527 44200
rect 6903 44252 6959 44254
rect 6903 44200 6905 44252
rect 6905 44200 6957 44252
rect 6957 44200 6959 44252
rect 7285 44214 7287 44266
rect 7287 44214 7339 44266
rect 7339 44214 7341 44266
rect 7285 44212 7341 44214
rect 7681 44266 7737 44268
rect 7681 44214 7683 44266
rect 7683 44214 7735 44266
rect 7735 44214 7737 44266
rect 7681 44212 7737 44214
rect 6903 44198 6959 44200
rect 6046 43894 6102 43896
rect 6046 43842 6048 43894
rect 6048 43842 6100 43894
rect 6100 43842 6102 43894
rect 6046 43840 6102 43842
rect 6471 43894 6527 43896
rect 6471 43842 6473 43894
rect 6473 43842 6525 43894
rect 6525 43842 6527 43894
rect 6471 43840 6527 43842
rect 6903 43894 6959 43896
rect 6903 43842 6905 43894
rect 6905 43842 6957 43894
rect 6957 43842 6959 43894
rect 6903 43840 6959 43842
rect 7285 43871 7341 43873
rect 7285 43819 7287 43871
rect 7287 43819 7339 43871
rect 7339 43819 7341 43871
rect 7285 43817 7341 43819
rect 7681 43871 7737 43873
rect 7681 43819 7683 43871
rect 7683 43819 7735 43871
rect 7735 43819 7737 43871
rect 7681 43817 7737 43819
rect 6046 43520 6102 43522
rect 6046 43468 6048 43520
rect 6048 43468 6100 43520
rect 6100 43468 6102 43520
rect 7285 43476 7341 43478
rect 6046 43466 6102 43468
rect 6471 43462 6527 43464
rect 6471 43410 6473 43462
rect 6473 43410 6525 43462
rect 6525 43410 6527 43462
rect 6471 43408 6527 43410
rect 6903 43462 6959 43464
rect 6903 43410 6905 43462
rect 6905 43410 6957 43462
rect 6957 43410 6959 43462
rect 7285 43424 7287 43476
rect 7287 43424 7339 43476
rect 7339 43424 7341 43476
rect 7285 43422 7341 43424
rect 7681 43476 7737 43478
rect 7681 43424 7683 43476
rect 7683 43424 7735 43476
rect 7735 43424 7737 43476
rect 7681 43422 7737 43424
rect 6903 43408 6959 43410
rect 6046 43104 6102 43106
rect 6046 43052 6048 43104
rect 6048 43052 6100 43104
rect 6100 43052 6102 43104
rect 6046 43050 6102 43052
rect 6471 43104 6527 43106
rect 6471 43052 6473 43104
rect 6473 43052 6525 43104
rect 6525 43052 6527 43104
rect 6471 43050 6527 43052
rect 6903 43104 6959 43106
rect 6903 43052 6905 43104
rect 6905 43052 6957 43104
rect 6957 43052 6959 43104
rect 6903 43050 6959 43052
rect 7285 43081 7341 43083
rect 7285 43029 7287 43081
rect 7287 43029 7339 43081
rect 7339 43029 7341 43081
rect 7285 43027 7341 43029
rect 7681 43081 7737 43083
rect 7681 43029 7683 43081
rect 7683 43029 7735 43081
rect 7735 43029 7737 43081
rect 7681 43027 7737 43029
rect 6046 42730 6102 42732
rect 6046 42678 6048 42730
rect 6048 42678 6100 42730
rect 6100 42678 6102 42730
rect 7285 42686 7341 42688
rect 6046 42676 6102 42678
rect 6471 42672 6527 42674
rect 6471 42620 6473 42672
rect 6473 42620 6525 42672
rect 6525 42620 6527 42672
rect 6471 42618 6527 42620
rect 6903 42672 6959 42674
rect 6903 42620 6905 42672
rect 6905 42620 6957 42672
rect 6957 42620 6959 42672
rect 7285 42634 7287 42686
rect 7287 42634 7339 42686
rect 7339 42634 7341 42686
rect 7285 42632 7341 42634
rect 7681 42686 7737 42688
rect 7681 42634 7683 42686
rect 7683 42634 7735 42686
rect 7735 42634 7737 42686
rect 7681 42632 7737 42634
rect 6903 42618 6959 42620
rect 6046 42314 6102 42316
rect 6046 42262 6048 42314
rect 6048 42262 6100 42314
rect 6100 42262 6102 42314
rect 6046 42260 6102 42262
rect 6471 42314 6527 42316
rect 6471 42262 6473 42314
rect 6473 42262 6525 42314
rect 6525 42262 6527 42314
rect 6471 42260 6527 42262
rect 6903 42314 6959 42316
rect 6903 42262 6905 42314
rect 6905 42262 6957 42314
rect 6957 42262 6959 42314
rect 6903 42260 6959 42262
rect 7285 42291 7341 42293
rect 7285 42239 7287 42291
rect 7287 42239 7339 42291
rect 7339 42239 7341 42291
rect 7285 42237 7341 42239
rect 7681 42291 7737 42293
rect 7681 42239 7683 42291
rect 7683 42239 7735 42291
rect 7735 42239 7737 42291
rect 7681 42237 7737 42239
rect 6046 41940 6102 41942
rect 6046 41888 6048 41940
rect 6048 41888 6100 41940
rect 6100 41888 6102 41940
rect 7285 41896 7341 41898
rect 6046 41886 6102 41888
rect 6471 41882 6527 41884
rect 6471 41830 6473 41882
rect 6473 41830 6525 41882
rect 6525 41830 6527 41882
rect 6471 41828 6527 41830
rect 6903 41882 6959 41884
rect 6903 41830 6905 41882
rect 6905 41830 6957 41882
rect 6957 41830 6959 41882
rect 7285 41844 7287 41896
rect 7287 41844 7339 41896
rect 7339 41844 7341 41896
rect 7285 41842 7341 41844
rect 7681 41896 7737 41898
rect 7681 41844 7683 41896
rect 7683 41844 7735 41896
rect 7735 41844 7737 41896
rect 7681 41842 7737 41844
rect 6903 41828 6959 41830
rect 6046 41524 6102 41526
rect 6046 41472 6048 41524
rect 6048 41472 6100 41524
rect 6100 41472 6102 41524
rect 6046 41470 6102 41472
rect 6471 41524 6527 41526
rect 6471 41472 6473 41524
rect 6473 41472 6525 41524
rect 6525 41472 6527 41524
rect 6471 41470 6527 41472
rect 6903 41524 6959 41526
rect 6903 41472 6905 41524
rect 6905 41472 6957 41524
rect 6957 41472 6959 41524
rect 6903 41470 6959 41472
rect 7285 41501 7341 41503
rect 7285 41449 7287 41501
rect 7287 41449 7339 41501
rect 7339 41449 7341 41501
rect 7285 41447 7341 41449
rect 7681 41501 7737 41503
rect 7681 41449 7683 41501
rect 7683 41449 7735 41501
rect 7735 41449 7737 41501
rect 7681 41447 7737 41449
rect 6046 41150 6102 41152
rect 6046 41098 6048 41150
rect 6048 41098 6100 41150
rect 6100 41098 6102 41150
rect 7285 41106 7341 41108
rect 6046 41096 6102 41098
rect 6471 41092 6527 41094
rect 6471 41040 6473 41092
rect 6473 41040 6525 41092
rect 6525 41040 6527 41092
rect 6471 41038 6527 41040
rect 6903 41092 6959 41094
rect 6903 41040 6905 41092
rect 6905 41040 6957 41092
rect 6957 41040 6959 41092
rect 7285 41054 7287 41106
rect 7287 41054 7339 41106
rect 7339 41054 7341 41106
rect 7285 41052 7341 41054
rect 7681 41106 7737 41108
rect 7681 41054 7683 41106
rect 7683 41054 7735 41106
rect 7735 41054 7737 41106
rect 7681 41052 7737 41054
rect 6903 41038 6959 41040
rect 6046 40734 6102 40736
rect 6046 40682 6048 40734
rect 6048 40682 6100 40734
rect 6100 40682 6102 40734
rect 6046 40680 6102 40682
rect 6471 40734 6527 40736
rect 6471 40682 6473 40734
rect 6473 40682 6525 40734
rect 6525 40682 6527 40734
rect 6471 40680 6527 40682
rect 6903 40734 6959 40736
rect 6903 40682 6905 40734
rect 6905 40682 6957 40734
rect 6957 40682 6959 40734
rect 6903 40680 6959 40682
rect 7285 40711 7341 40713
rect 7285 40659 7287 40711
rect 7287 40659 7339 40711
rect 7339 40659 7341 40711
rect 7285 40657 7341 40659
rect 7681 40711 7737 40713
rect 7681 40659 7683 40711
rect 7683 40659 7735 40711
rect 7735 40659 7737 40711
rect 7681 40657 7737 40659
rect 6046 40360 6102 40362
rect 6046 40308 6048 40360
rect 6048 40308 6100 40360
rect 6100 40308 6102 40360
rect 7285 40316 7341 40318
rect 6046 40306 6102 40308
rect 6471 40302 6527 40304
rect 6471 40250 6473 40302
rect 6473 40250 6525 40302
rect 6525 40250 6527 40302
rect 6471 40248 6527 40250
rect 6903 40302 6959 40304
rect 6903 40250 6905 40302
rect 6905 40250 6957 40302
rect 6957 40250 6959 40302
rect 7285 40264 7287 40316
rect 7287 40264 7339 40316
rect 7339 40264 7341 40316
rect 7285 40262 7341 40264
rect 7681 40316 7737 40318
rect 7681 40264 7683 40316
rect 7683 40264 7735 40316
rect 7735 40264 7737 40316
rect 7681 40262 7737 40264
rect 6903 40248 6959 40250
rect 6046 39944 6102 39946
rect 6046 39892 6048 39944
rect 6048 39892 6100 39944
rect 6100 39892 6102 39944
rect 6046 39890 6102 39892
rect 6471 39944 6527 39946
rect 6471 39892 6473 39944
rect 6473 39892 6525 39944
rect 6525 39892 6527 39944
rect 6471 39890 6527 39892
rect 6903 39944 6959 39946
rect 6903 39892 6905 39944
rect 6905 39892 6957 39944
rect 6957 39892 6959 39944
rect 6903 39890 6959 39892
rect 7285 39921 7341 39923
rect 7285 39869 7287 39921
rect 7287 39869 7339 39921
rect 7339 39869 7341 39921
rect 7285 39867 7341 39869
rect 7681 39921 7737 39923
rect 7681 39869 7683 39921
rect 7683 39869 7735 39921
rect 7735 39869 7737 39921
rect 7681 39867 7737 39869
rect 6046 39570 6102 39572
rect 6046 39518 6048 39570
rect 6048 39518 6100 39570
rect 6100 39518 6102 39570
rect 7285 39526 7341 39528
rect 6046 39516 6102 39518
rect 6471 39512 6527 39514
rect 6471 39460 6473 39512
rect 6473 39460 6525 39512
rect 6525 39460 6527 39512
rect 6471 39458 6527 39460
rect 6903 39512 6959 39514
rect 6903 39460 6905 39512
rect 6905 39460 6957 39512
rect 6957 39460 6959 39512
rect 7285 39474 7287 39526
rect 7287 39474 7339 39526
rect 7339 39474 7341 39526
rect 7285 39472 7341 39474
rect 7681 39526 7737 39528
rect 7681 39474 7683 39526
rect 7683 39474 7735 39526
rect 7735 39474 7737 39526
rect 7681 39472 7737 39474
rect 6903 39458 6959 39460
rect 6046 39154 6102 39156
rect 6046 39102 6048 39154
rect 6048 39102 6100 39154
rect 6100 39102 6102 39154
rect 6046 39100 6102 39102
rect 6471 39154 6527 39156
rect 6471 39102 6473 39154
rect 6473 39102 6525 39154
rect 6525 39102 6527 39154
rect 6471 39100 6527 39102
rect 6903 39154 6959 39156
rect 6903 39102 6905 39154
rect 6905 39102 6957 39154
rect 6957 39102 6959 39154
rect 6903 39100 6959 39102
rect 7285 39131 7341 39133
rect 7285 39079 7287 39131
rect 7287 39079 7339 39131
rect 7339 39079 7341 39131
rect 7285 39077 7341 39079
rect 7681 39131 7737 39133
rect 7681 39079 7683 39131
rect 7683 39079 7735 39131
rect 7735 39079 7737 39131
rect 7681 39077 7737 39079
rect 6046 38780 6102 38782
rect 6046 38728 6048 38780
rect 6048 38728 6100 38780
rect 6100 38728 6102 38780
rect 7285 38736 7341 38738
rect 6046 38726 6102 38728
rect 6471 38722 6527 38724
rect 6471 38670 6473 38722
rect 6473 38670 6525 38722
rect 6525 38670 6527 38722
rect 6471 38668 6527 38670
rect 6903 38722 6959 38724
rect 6903 38670 6905 38722
rect 6905 38670 6957 38722
rect 6957 38670 6959 38722
rect 7285 38684 7287 38736
rect 7287 38684 7339 38736
rect 7339 38684 7341 38736
rect 7285 38682 7341 38684
rect 7681 38736 7737 38738
rect 7681 38684 7683 38736
rect 7683 38684 7735 38736
rect 7735 38684 7737 38736
rect 7681 38682 7737 38684
rect 6903 38668 6959 38670
rect 6046 38364 6102 38366
rect 6046 38312 6048 38364
rect 6048 38312 6100 38364
rect 6100 38312 6102 38364
rect 6046 38310 6102 38312
rect 6471 38364 6527 38366
rect 6471 38312 6473 38364
rect 6473 38312 6525 38364
rect 6525 38312 6527 38364
rect 6471 38310 6527 38312
rect 6903 38364 6959 38366
rect 6903 38312 6905 38364
rect 6905 38312 6957 38364
rect 6957 38312 6959 38364
rect 6903 38310 6959 38312
rect 7285 38341 7341 38343
rect 7285 38289 7287 38341
rect 7287 38289 7339 38341
rect 7339 38289 7341 38341
rect 7285 38287 7341 38289
rect 7681 38341 7737 38343
rect 7681 38289 7683 38341
rect 7683 38289 7735 38341
rect 7735 38289 7737 38341
rect 7681 38287 7737 38289
rect 6046 37990 6102 37992
rect 6046 37938 6048 37990
rect 6048 37938 6100 37990
rect 6100 37938 6102 37990
rect 7285 37946 7341 37948
rect 6046 37936 6102 37938
rect 6471 37932 6527 37934
rect 6471 37880 6473 37932
rect 6473 37880 6525 37932
rect 6525 37880 6527 37932
rect 6471 37878 6527 37880
rect 6903 37932 6959 37934
rect 6903 37880 6905 37932
rect 6905 37880 6957 37932
rect 6957 37880 6959 37932
rect 7285 37894 7287 37946
rect 7287 37894 7339 37946
rect 7339 37894 7341 37946
rect 7285 37892 7341 37894
rect 7681 37946 7737 37948
rect 7681 37894 7683 37946
rect 7683 37894 7735 37946
rect 7735 37894 7737 37946
rect 7681 37892 7737 37894
rect 6903 37878 6959 37880
rect 6046 37574 6102 37576
rect 6046 37522 6048 37574
rect 6048 37522 6100 37574
rect 6100 37522 6102 37574
rect 6046 37520 6102 37522
rect 6471 37574 6527 37576
rect 6471 37522 6473 37574
rect 6473 37522 6525 37574
rect 6525 37522 6527 37574
rect 6471 37520 6527 37522
rect 6903 37574 6959 37576
rect 6903 37522 6905 37574
rect 6905 37522 6957 37574
rect 6957 37522 6959 37574
rect 6903 37520 6959 37522
rect 7285 37551 7341 37553
rect 7285 37499 7287 37551
rect 7287 37499 7339 37551
rect 7339 37499 7341 37551
rect 7285 37497 7341 37499
rect 7681 37551 7737 37553
rect 7681 37499 7683 37551
rect 7683 37499 7735 37551
rect 7735 37499 7737 37551
rect 7681 37497 7737 37499
rect 6046 37200 6102 37202
rect 6046 37148 6048 37200
rect 6048 37148 6100 37200
rect 6100 37148 6102 37200
rect 7285 37156 7341 37158
rect 6046 37146 6102 37148
rect 6471 37142 6527 37144
rect 6471 37090 6473 37142
rect 6473 37090 6525 37142
rect 6525 37090 6527 37142
rect 6471 37088 6527 37090
rect 6903 37142 6959 37144
rect 6903 37090 6905 37142
rect 6905 37090 6957 37142
rect 6957 37090 6959 37142
rect 7285 37104 7287 37156
rect 7287 37104 7339 37156
rect 7339 37104 7341 37156
rect 7285 37102 7341 37104
rect 7681 37156 7737 37158
rect 7681 37104 7683 37156
rect 7683 37104 7735 37156
rect 7735 37104 7737 37156
rect 7681 37102 7737 37104
rect 6903 37088 6959 37090
rect 6046 36784 6102 36786
rect 6046 36732 6048 36784
rect 6048 36732 6100 36784
rect 6100 36732 6102 36784
rect 6046 36730 6102 36732
rect 6471 36784 6527 36786
rect 6471 36732 6473 36784
rect 6473 36732 6525 36784
rect 6525 36732 6527 36784
rect 6471 36730 6527 36732
rect 6903 36784 6959 36786
rect 6903 36732 6905 36784
rect 6905 36732 6957 36784
rect 6957 36732 6959 36784
rect 6903 36730 6959 36732
rect 7285 36761 7341 36763
rect 7285 36709 7287 36761
rect 7287 36709 7339 36761
rect 7339 36709 7341 36761
rect 7285 36707 7341 36709
rect 7681 36761 7737 36763
rect 7681 36709 7683 36761
rect 7683 36709 7735 36761
rect 7735 36709 7737 36761
rect 7681 36707 7737 36709
rect 6046 36410 6102 36412
rect 6046 36358 6048 36410
rect 6048 36358 6100 36410
rect 6100 36358 6102 36410
rect 7285 36366 7341 36368
rect 6046 36356 6102 36358
rect 6471 36352 6527 36354
rect 6471 36300 6473 36352
rect 6473 36300 6525 36352
rect 6525 36300 6527 36352
rect 6471 36298 6527 36300
rect 6903 36352 6959 36354
rect 6903 36300 6905 36352
rect 6905 36300 6957 36352
rect 6957 36300 6959 36352
rect 7285 36314 7287 36366
rect 7287 36314 7339 36366
rect 7339 36314 7341 36366
rect 7285 36312 7341 36314
rect 7681 36366 7737 36368
rect 7681 36314 7683 36366
rect 7683 36314 7735 36366
rect 7735 36314 7737 36366
rect 7681 36312 7737 36314
rect 6903 36298 6959 36300
rect 6046 35994 6102 35996
rect 6046 35942 6048 35994
rect 6048 35942 6100 35994
rect 6100 35942 6102 35994
rect 6046 35940 6102 35942
rect 6471 35994 6527 35996
rect 6471 35942 6473 35994
rect 6473 35942 6525 35994
rect 6525 35942 6527 35994
rect 6471 35940 6527 35942
rect 6903 35994 6959 35996
rect 6903 35942 6905 35994
rect 6905 35942 6957 35994
rect 6957 35942 6959 35994
rect 6903 35940 6959 35942
rect 7285 35971 7341 35973
rect 7285 35919 7287 35971
rect 7287 35919 7339 35971
rect 7339 35919 7341 35971
rect 7285 35917 7341 35919
rect 7681 35971 7737 35973
rect 7681 35919 7683 35971
rect 7683 35919 7735 35971
rect 7735 35919 7737 35971
rect 7681 35917 7737 35919
rect 6046 35620 6102 35622
rect 6046 35568 6048 35620
rect 6048 35568 6100 35620
rect 6100 35568 6102 35620
rect 7285 35576 7341 35578
rect 6046 35566 6102 35568
rect 6471 35562 6527 35564
rect 6471 35510 6473 35562
rect 6473 35510 6525 35562
rect 6525 35510 6527 35562
rect 6471 35508 6527 35510
rect 6903 35562 6959 35564
rect 6903 35510 6905 35562
rect 6905 35510 6957 35562
rect 6957 35510 6959 35562
rect 7285 35524 7287 35576
rect 7287 35524 7339 35576
rect 7339 35524 7341 35576
rect 7285 35522 7341 35524
rect 7681 35576 7737 35578
rect 7681 35524 7683 35576
rect 7683 35524 7735 35576
rect 7735 35524 7737 35576
rect 7681 35522 7737 35524
rect 6903 35508 6959 35510
rect 6046 35204 6102 35206
rect 6046 35152 6048 35204
rect 6048 35152 6100 35204
rect 6100 35152 6102 35204
rect 6046 35150 6102 35152
rect 6471 35204 6527 35206
rect 6471 35152 6473 35204
rect 6473 35152 6525 35204
rect 6525 35152 6527 35204
rect 6471 35150 6527 35152
rect 6903 35204 6959 35206
rect 6903 35152 6905 35204
rect 6905 35152 6957 35204
rect 6957 35152 6959 35204
rect 6903 35150 6959 35152
rect 7285 35181 7341 35183
rect 7285 35129 7287 35181
rect 7287 35129 7339 35181
rect 7339 35129 7341 35181
rect 7285 35127 7341 35129
rect 7681 35181 7737 35183
rect 7681 35129 7683 35181
rect 7683 35129 7735 35181
rect 7735 35129 7737 35181
rect 7681 35127 7737 35129
rect 6046 34830 6102 34832
rect 6046 34778 6048 34830
rect 6048 34778 6100 34830
rect 6100 34778 6102 34830
rect 7285 34786 7341 34788
rect 6046 34776 6102 34778
rect 6471 34772 6527 34774
rect 6471 34720 6473 34772
rect 6473 34720 6525 34772
rect 6525 34720 6527 34772
rect 6471 34718 6527 34720
rect 6903 34772 6959 34774
rect 6903 34720 6905 34772
rect 6905 34720 6957 34772
rect 6957 34720 6959 34772
rect 7285 34734 7287 34786
rect 7287 34734 7339 34786
rect 7339 34734 7341 34786
rect 7285 34732 7341 34734
rect 7681 34786 7737 34788
rect 7681 34734 7683 34786
rect 7683 34734 7735 34786
rect 7735 34734 7737 34786
rect 7681 34732 7737 34734
rect 6903 34718 6959 34720
rect 6046 34414 6102 34416
rect 6046 34362 6048 34414
rect 6048 34362 6100 34414
rect 6100 34362 6102 34414
rect 6046 34360 6102 34362
rect 6471 34414 6527 34416
rect 6471 34362 6473 34414
rect 6473 34362 6525 34414
rect 6525 34362 6527 34414
rect 6471 34360 6527 34362
rect 6903 34414 6959 34416
rect 6903 34362 6905 34414
rect 6905 34362 6957 34414
rect 6957 34362 6959 34414
rect 6903 34360 6959 34362
rect 7285 34391 7341 34393
rect 7285 34339 7287 34391
rect 7287 34339 7339 34391
rect 7339 34339 7341 34391
rect 7285 34337 7341 34339
rect 7681 34391 7737 34393
rect 7681 34339 7683 34391
rect 7683 34339 7735 34391
rect 7735 34339 7737 34391
rect 7681 34337 7737 34339
rect 6046 34040 6102 34042
rect 6046 33988 6048 34040
rect 6048 33988 6100 34040
rect 6100 33988 6102 34040
rect 7285 33996 7341 33998
rect 6046 33986 6102 33988
rect 6471 33982 6527 33984
rect 6471 33930 6473 33982
rect 6473 33930 6525 33982
rect 6525 33930 6527 33982
rect 6471 33928 6527 33930
rect 6903 33982 6959 33984
rect 6903 33930 6905 33982
rect 6905 33930 6957 33982
rect 6957 33930 6959 33982
rect 7285 33944 7287 33996
rect 7287 33944 7339 33996
rect 7339 33944 7341 33996
rect 7285 33942 7341 33944
rect 7681 33996 7737 33998
rect 7681 33944 7683 33996
rect 7683 33944 7735 33996
rect 7735 33944 7737 33996
rect 7681 33942 7737 33944
rect 6903 33928 6959 33930
rect 6046 33624 6102 33626
rect 6046 33572 6048 33624
rect 6048 33572 6100 33624
rect 6100 33572 6102 33624
rect 6046 33570 6102 33572
rect 6471 33624 6527 33626
rect 6471 33572 6473 33624
rect 6473 33572 6525 33624
rect 6525 33572 6527 33624
rect 6471 33570 6527 33572
rect 6903 33624 6959 33626
rect 6903 33572 6905 33624
rect 6905 33572 6957 33624
rect 6957 33572 6959 33624
rect 6903 33570 6959 33572
rect 7285 33601 7341 33603
rect 7285 33549 7287 33601
rect 7287 33549 7339 33601
rect 7339 33549 7341 33601
rect 7285 33547 7341 33549
rect 7681 33601 7737 33603
rect 7681 33549 7683 33601
rect 7683 33549 7735 33601
rect 7735 33549 7737 33601
rect 7681 33547 7737 33549
rect 6046 33250 6102 33252
rect 6046 33198 6048 33250
rect 6048 33198 6100 33250
rect 6100 33198 6102 33250
rect 7285 33206 7341 33208
rect 6046 33196 6102 33198
rect 6471 33192 6527 33194
rect 6471 33140 6473 33192
rect 6473 33140 6525 33192
rect 6525 33140 6527 33192
rect 6471 33138 6527 33140
rect 6903 33192 6959 33194
rect 6903 33140 6905 33192
rect 6905 33140 6957 33192
rect 6957 33140 6959 33192
rect 7285 33154 7287 33206
rect 7287 33154 7339 33206
rect 7339 33154 7341 33206
rect 7285 33152 7341 33154
rect 7681 33206 7737 33208
rect 7681 33154 7683 33206
rect 7683 33154 7735 33206
rect 7735 33154 7737 33206
rect 7681 33152 7737 33154
rect 6903 33138 6959 33140
rect 6046 32834 6102 32836
rect 6046 32782 6048 32834
rect 6048 32782 6100 32834
rect 6100 32782 6102 32834
rect 6046 32780 6102 32782
rect 6471 32834 6527 32836
rect 6471 32782 6473 32834
rect 6473 32782 6525 32834
rect 6525 32782 6527 32834
rect 6471 32780 6527 32782
rect 6903 32834 6959 32836
rect 6903 32782 6905 32834
rect 6905 32782 6957 32834
rect 6957 32782 6959 32834
rect 6903 32780 6959 32782
rect 7285 32811 7341 32813
rect 7285 32759 7287 32811
rect 7287 32759 7339 32811
rect 7339 32759 7341 32811
rect 7285 32757 7341 32759
rect 7681 32811 7737 32813
rect 7681 32759 7683 32811
rect 7683 32759 7735 32811
rect 7735 32759 7737 32811
rect 7681 32757 7737 32759
rect 6046 32460 6102 32462
rect 6046 32408 6048 32460
rect 6048 32408 6100 32460
rect 6100 32408 6102 32460
rect 7285 32416 7341 32418
rect 6046 32406 6102 32408
rect 6471 32402 6527 32404
rect 6471 32350 6473 32402
rect 6473 32350 6525 32402
rect 6525 32350 6527 32402
rect 6471 32348 6527 32350
rect 6903 32402 6959 32404
rect 6903 32350 6905 32402
rect 6905 32350 6957 32402
rect 6957 32350 6959 32402
rect 7285 32364 7287 32416
rect 7287 32364 7339 32416
rect 7339 32364 7341 32416
rect 7285 32362 7341 32364
rect 7681 32416 7737 32418
rect 7681 32364 7683 32416
rect 7683 32364 7735 32416
rect 7735 32364 7737 32416
rect 7681 32362 7737 32364
rect 6903 32348 6959 32350
rect 6046 32044 6102 32046
rect 6046 31992 6048 32044
rect 6048 31992 6100 32044
rect 6100 31992 6102 32044
rect 6046 31990 6102 31992
rect 6471 32044 6527 32046
rect 6471 31992 6473 32044
rect 6473 31992 6525 32044
rect 6525 31992 6527 32044
rect 6471 31990 6527 31992
rect 6903 32044 6959 32046
rect 6903 31992 6905 32044
rect 6905 31992 6957 32044
rect 6957 31992 6959 32044
rect 6903 31990 6959 31992
rect 7285 32021 7341 32023
rect 7285 31969 7287 32021
rect 7287 31969 7339 32021
rect 7339 31969 7341 32021
rect 7285 31967 7341 31969
rect 7681 32021 7737 32023
rect 7681 31969 7683 32021
rect 7683 31969 7735 32021
rect 7735 31969 7737 32021
rect 7681 31967 7737 31969
rect 6046 31670 6102 31672
rect 6046 31618 6048 31670
rect 6048 31618 6100 31670
rect 6100 31618 6102 31670
rect 7285 31626 7341 31628
rect 6046 31616 6102 31618
rect 6471 31612 6527 31614
rect 6471 31560 6473 31612
rect 6473 31560 6525 31612
rect 6525 31560 6527 31612
rect 6471 31558 6527 31560
rect 6903 31612 6959 31614
rect 6903 31560 6905 31612
rect 6905 31560 6957 31612
rect 6957 31560 6959 31612
rect 7285 31574 7287 31626
rect 7287 31574 7339 31626
rect 7339 31574 7341 31626
rect 7285 31572 7341 31574
rect 7681 31626 7737 31628
rect 7681 31574 7683 31626
rect 7683 31574 7735 31626
rect 7735 31574 7737 31626
rect 7681 31572 7737 31574
rect 6903 31558 6959 31560
rect 6046 31254 6102 31256
rect 6046 31202 6048 31254
rect 6048 31202 6100 31254
rect 6100 31202 6102 31254
rect 6046 31200 6102 31202
rect 6471 31254 6527 31256
rect 6471 31202 6473 31254
rect 6473 31202 6525 31254
rect 6525 31202 6527 31254
rect 6471 31200 6527 31202
rect 6903 31254 6959 31256
rect 6903 31202 6905 31254
rect 6905 31202 6957 31254
rect 6957 31202 6959 31254
rect 6903 31200 6959 31202
rect 7285 31231 7341 31233
rect 7285 31179 7287 31231
rect 7287 31179 7339 31231
rect 7339 31179 7341 31231
rect 7285 31177 7341 31179
rect 7681 31231 7737 31233
rect 7681 31179 7683 31231
rect 7683 31179 7735 31231
rect 7735 31179 7737 31231
rect 7681 31177 7737 31179
rect 6046 30880 6102 30882
rect 6046 30828 6048 30880
rect 6048 30828 6100 30880
rect 6100 30828 6102 30880
rect 7285 30836 7341 30838
rect 6046 30826 6102 30828
rect 6471 30822 6527 30824
rect 6471 30770 6473 30822
rect 6473 30770 6525 30822
rect 6525 30770 6527 30822
rect 6471 30768 6527 30770
rect 6903 30822 6959 30824
rect 6903 30770 6905 30822
rect 6905 30770 6957 30822
rect 6957 30770 6959 30822
rect 7285 30784 7287 30836
rect 7287 30784 7339 30836
rect 7339 30784 7341 30836
rect 7285 30782 7341 30784
rect 7681 30836 7737 30838
rect 7681 30784 7683 30836
rect 7683 30784 7735 30836
rect 7735 30784 7737 30836
rect 7681 30782 7737 30784
rect 6903 30768 6959 30770
rect 6046 30464 6102 30466
rect 6046 30412 6048 30464
rect 6048 30412 6100 30464
rect 6100 30412 6102 30464
rect 6046 30410 6102 30412
rect 6471 30464 6527 30466
rect 6471 30412 6473 30464
rect 6473 30412 6525 30464
rect 6525 30412 6527 30464
rect 6471 30410 6527 30412
rect 6903 30464 6959 30466
rect 6903 30412 6905 30464
rect 6905 30412 6957 30464
rect 6957 30412 6959 30464
rect 6903 30410 6959 30412
rect 7285 30441 7341 30443
rect 7285 30389 7287 30441
rect 7287 30389 7339 30441
rect 7339 30389 7341 30441
rect 7285 30387 7341 30389
rect 7681 30441 7737 30443
rect 7681 30389 7683 30441
rect 7683 30389 7735 30441
rect 7735 30389 7737 30441
rect 7681 30387 7737 30389
rect 6046 30090 6102 30092
rect 6046 30038 6048 30090
rect 6048 30038 6100 30090
rect 6100 30038 6102 30090
rect 7285 30046 7341 30048
rect 6046 30036 6102 30038
rect 6471 30032 6527 30034
rect 6471 29980 6473 30032
rect 6473 29980 6525 30032
rect 6525 29980 6527 30032
rect 6471 29978 6527 29980
rect 6903 30032 6959 30034
rect 6903 29980 6905 30032
rect 6905 29980 6957 30032
rect 6957 29980 6959 30032
rect 7285 29994 7287 30046
rect 7287 29994 7339 30046
rect 7339 29994 7341 30046
rect 7285 29992 7341 29994
rect 7681 30046 7737 30048
rect 7681 29994 7683 30046
rect 7683 29994 7735 30046
rect 7735 29994 7737 30046
rect 7681 29992 7737 29994
rect 6903 29978 6959 29980
rect 6046 29674 6102 29676
rect 6046 29622 6048 29674
rect 6048 29622 6100 29674
rect 6100 29622 6102 29674
rect 6046 29620 6102 29622
rect 6471 29674 6527 29676
rect 6471 29622 6473 29674
rect 6473 29622 6525 29674
rect 6525 29622 6527 29674
rect 6471 29620 6527 29622
rect 6903 29674 6959 29676
rect 6903 29622 6905 29674
rect 6905 29622 6957 29674
rect 6957 29622 6959 29674
rect 6903 29620 6959 29622
rect 7285 29651 7341 29653
rect 7285 29599 7287 29651
rect 7287 29599 7339 29651
rect 7339 29599 7341 29651
rect 7285 29597 7341 29599
rect 7681 29651 7737 29653
rect 7681 29599 7683 29651
rect 7683 29599 7735 29651
rect 7735 29599 7737 29651
rect 7681 29597 7737 29599
rect 6046 29300 6102 29302
rect 6046 29248 6048 29300
rect 6048 29248 6100 29300
rect 6100 29248 6102 29300
rect 7285 29256 7341 29258
rect 6046 29246 6102 29248
rect 6471 29242 6527 29244
rect 6471 29190 6473 29242
rect 6473 29190 6525 29242
rect 6525 29190 6527 29242
rect 6471 29188 6527 29190
rect 6903 29242 6959 29244
rect 6903 29190 6905 29242
rect 6905 29190 6957 29242
rect 6957 29190 6959 29242
rect 7285 29204 7287 29256
rect 7287 29204 7339 29256
rect 7339 29204 7341 29256
rect 7285 29202 7341 29204
rect 7681 29256 7737 29258
rect 7681 29204 7683 29256
rect 7683 29204 7735 29256
rect 7735 29204 7737 29256
rect 7681 29202 7737 29204
rect 6903 29188 6959 29190
rect 6046 28884 6102 28886
rect 6046 28832 6048 28884
rect 6048 28832 6100 28884
rect 6100 28832 6102 28884
rect 6046 28830 6102 28832
rect 6471 28884 6527 28886
rect 6471 28832 6473 28884
rect 6473 28832 6525 28884
rect 6525 28832 6527 28884
rect 6471 28830 6527 28832
rect 6903 28884 6959 28886
rect 6903 28832 6905 28884
rect 6905 28832 6957 28884
rect 6957 28832 6959 28884
rect 6903 28830 6959 28832
rect 7285 28861 7341 28863
rect 7285 28809 7287 28861
rect 7287 28809 7339 28861
rect 7339 28809 7341 28861
rect 7285 28807 7341 28809
rect 7681 28861 7737 28863
rect 7681 28809 7683 28861
rect 7683 28809 7735 28861
rect 7735 28809 7737 28861
rect 7681 28807 7737 28809
rect 6046 28510 6102 28512
rect 6046 28458 6048 28510
rect 6048 28458 6100 28510
rect 6100 28458 6102 28510
rect 7285 28466 7341 28468
rect 6046 28456 6102 28458
rect 6471 28452 6527 28454
rect 6471 28400 6473 28452
rect 6473 28400 6525 28452
rect 6525 28400 6527 28452
rect 6471 28398 6527 28400
rect 6903 28452 6959 28454
rect 6903 28400 6905 28452
rect 6905 28400 6957 28452
rect 6957 28400 6959 28452
rect 7285 28414 7287 28466
rect 7287 28414 7339 28466
rect 7339 28414 7341 28466
rect 7285 28412 7341 28414
rect 7681 28466 7737 28468
rect 7681 28414 7683 28466
rect 7683 28414 7735 28466
rect 7735 28414 7737 28466
rect 7681 28412 7737 28414
rect 6903 28398 6959 28400
rect 6046 28094 6102 28096
rect 6046 28042 6048 28094
rect 6048 28042 6100 28094
rect 6100 28042 6102 28094
rect 6046 28040 6102 28042
rect 6471 28094 6527 28096
rect 6471 28042 6473 28094
rect 6473 28042 6525 28094
rect 6525 28042 6527 28094
rect 6471 28040 6527 28042
rect 6903 28094 6959 28096
rect 6903 28042 6905 28094
rect 6905 28042 6957 28094
rect 6957 28042 6959 28094
rect 6903 28040 6959 28042
rect 7285 28071 7341 28073
rect 7285 28019 7287 28071
rect 7287 28019 7339 28071
rect 7339 28019 7341 28071
rect 7285 28017 7341 28019
rect 7681 28071 7737 28073
rect 7681 28019 7683 28071
rect 7683 28019 7735 28071
rect 7735 28019 7737 28071
rect 7681 28017 7737 28019
rect 6046 27720 6102 27722
rect 6046 27668 6048 27720
rect 6048 27668 6100 27720
rect 6100 27668 6102 27720
rect 7285 27676 7341 27678
rect 6046 27666 6102 27668
rect 6471 27662 6527 27664
rect 6471 27610 6473 27662
rect 6473 27610 6525 27662
rect 6525 27610 6527 27662
rect 6471 27608 6527 27610
rect 6903 27662 6959 27664
rect 6903 27610 6905 27662
rect 6905 27610 6957 27662
rect 6957 27610 6959 27662
rect 7285 27624 7287 27676
rect 7287 27624 7339 27676
rect 7339 27624 7341 27676
rect 7285 27622 7341 27624
rect 7681 27676 7737 27678
rect 7681 27624 7683 27676
rect 7683 27624 7735 27676
rect 7735 27624 7737 27676
rect 7681 27622 7737 27624
rect 6903 27608 6959 27610
rect 6046 27304 6102 27306
rect 6046 27252 6048 27304
rect 6048 27252 6100 27304
rect 6100 27252 6102 27304
rect 6046 27250 6102 27252
rect 6471 27304 6527 27306
rect 6471 27252 6473 27304
rect 6473 27252 6525 27304
rect 6525 27252 6527 27304
rect 6471 27250 6527 27252
rect 6903 27304 6959 27306
rect 6903 27252 6905 27304
rect 6905 27252 6957 27304
rect 6957 27252 6959 27304
rect 6903 27250 6959 27252
rect 7285 27281 7341 27283
rect 7285 27229 7287 27281
rect 7287 27229 7339 27281
rect 7339 27229 7341 27281
rect 7285 27227 7341 27229
rect 7681 27281 7737 27283
rect 7681 27229 7683 27281
rect 7683 27229 7735 27281
rect 7735 27229 7737 27281
rect 7681 27227 7737 27229
rect 6046 26930 6102 26932
rect 6046 26878 6048 26930
rect 6048 26878 6100 26930
rect 6100 26878 6102 26930
rect 7285 26886 7341 26888
rect 6046 26876 6102 26878
rect 6471 26872 6527 26874
rect 6471 26820 6473 26872
rect 6473 26820 6525 26872
rect 6525 26820 6527 26872
rect 6471 26818 6527 26820
rect 6903 26872 6959 26874
rect 6903 26820 6905 26872
rect 6905 26820 6957 26872
rect 6957 26820 6959 26872
rect 7285 26834 7287 26886
rect 7287 26834 7339 26886
rect 7339 26834 7341 26886
rect 7285 26832 7341 26834
rect 7681 26886 7737 26888
rect 7681 26834 7683 26886
rect 7683 26834 7735 26886
rect 7735 26834 7737 26886
rect 7681 26832 7737 26834
rect 6903 26818 6959 26820
rect 6046 26514 6102 26516
rect 6046 26462 6048 26514
rect 6048 26462 6100 26514
rect 6100 26462 6102 26514
rect 6046 26460 6102 26462
rect 6471 26514 6527 26516
rect 6471 26462 6473 26514
rect 6473 26462 6525 26514
rect 6525 26462 6527 26514
rect 6471 26460 6527 26462
rect 6903 26514 6959 26516
rect 6903 26462 6905 26514
rect 6905 26462 6957 26514
rect 6957 26462 6959 26514
rect 6903 26460 6959 26462
rect 7285 26491 7341 26493
rect 7285 26439 7287 26491
rect 7287 26439 7339 26491
rect 7339 26439 7341 26491
rect 7285 26437 7341 26439
rect 7681 26491 7737 26493
rect 7681 26439 7683 26491
rect 7683 26439 7735 26491
rect 7735 26439 7737 26491
rect 7681 26437 7737 26439
rect 6046 26140 6102 26142
rect 6046 26088 6048 26140
rect 6048 26088 6100 26140
rect 6100 26088 6102 26140
rect 7285 26096 7341 26098
rect 6046 26086 6102 26088
rect 6471 26082 6527 26084
rect 6471 26030 6473 26082
rect 6473 26030 6525 26082
rect 6525 26030 6527 26082
rect 6471 26028 6527 26030
rect 6903 26082 6959 26084
rect 6903 26030 6905 26082
rect 6905 26030 6957 26082
rect 6957 26030 6959 26082
rect 7285 26044 7287 26096
rect 7287 26044 7339 26096
rect 7339 26044 7341 26096
rect 7285 26042 7341 26044
rect 7681 26096 7737 26098
rect 7681 26044 7683 26096
rect 7683 26044 7735 26096
rect 7735 26044 7737 26096
rect 7681 26042 7737 26044
rect 6903 26028 6959 26030
rect 6046 25724 6102 25726
rect 6046 25672 6048 25724
rect 6048 25672 6100 25724
rect 6100 25672 6102 25724
rect 6046 25670 6102 25672
rect 6471 25724 6527 25726
rect 6471 25672 6473 25724
rect 6473 25672 6525 25724
rect 6525 25672 6527 25724
rect 6471 25670 6527 25672
rect 6903 25724 6959 25726
rect 6903 25672 6905 25724
rect 6905 25672 6957 25724
rect 6957 25672 6959 25724
rect 6903 25670 6959 25672
rect 7285 25701 7341 25703
rect 7285 25649 7287 25701
rect 7287 25649 7339 25701
rect 7339 25649 7341 25701
rect 7285 25647 7341 25649
rect 7681 25701 7737 25703
rect 7681 25649 7683 25701
rect 7683 25649 7735 25701
rect 7735 25649 7737 25701
rect 7681 25647 7737 25649
rect 6046 25350 6102 25352
rect 6046 25298 6048 25350
rect 6048 25298 6100 25350
rect 6100 25298 6102 25350
rect 7285 25306 7341 25308
rect 6046 25296 6102 25298
rect 6471 25292 6527 25294
rect 6471 25240 6473 25292
rect 6473 25240 6525 25292
rect 6525 25240 6527 25292
rect 6471 25238 6527 25240
rect 6903 25292 6959 25294
rect 6903 25240 6905 25292
rect 6905 25240 6957 25292
rect 6957 25240 6959 25292
rect 7285 25254 7287 25306
rect 7287 25254 7339 25306
rect 7339 25254 7341 25306
rect 7285 25252 7341 25254
rect 7681 25306 7737 25308
rect 7681 25254 7683 25306
rect 7683 25254 7735 25306
rect 7735 25254 7737 25306
rect 7681 25252 7737 25254
rect 6903 25238 6959 25240
rect 6046 24934 6102 24936
rect 6046 24882 6048 24934
rect 6048 24882 6100 24934
rect 6100 24882 6102 24934
rect 6046 24880 6102 24882
rect 6471 24934 6527 24936
rect 6471 24882 6473 24934
rect 6473 24882 6525 24934
rect 6525 24882 6527 24934
rect 6471 24880 6527 24882
rect 6903 24934 6959 24936
rect 6903 24882 6905 24934
rect 6905 24882 6957 24934
rect 6957 24882 6959 24934
rect 6903 24880 6959 24882
rect 7285 24911 7341 24913
rect 7285 24859 7287 24911
rect 7287 24859 7339 24911
rect 7339 24859 7341 24911
rect 7285 24857 7341 24859
rect 7681 24911 7737 24913
rect 7681 24859 7683 24911
rect 7683 24859 7735 24911
rect 7735 24859 7737 24911
rect 7681 24857 7737 24859
rect 6046 24560 6102 24562
rect 6046 24508 6048 24560
rect 6048 24508 6100 24560
rect 6100 24508 6102 24560
rect 7285 24516 7341 24518
rect 6046 24506 6102 24508
rect 6471 24502 6527 24504
rect 6471 24450 6473 24502
rect 6473 24450 6525 24502
rect 6525 24450 6527 24502
rect 6471 24448 6527 24450
rect 6903 24502 6959 24504
rect 6903 24450 6905 24502
rect 6905 24450 6957 24502
rect 6957 24450 6959 24502
rect 7285 24464 7287 24516
rect 7287 24464 7339 24516
rect 7339 24464 7341 24516
rect 7285 24462 7341 24464
rect 7681 24516 7737 24518
rect 7681 24464 7683 24516
rect 7683 24464 7735 24516
rect 7735 24464 7737 24516
rect 7681 24462 7737 24464
rect 6903 24448 6959 24450
rect 6046 24144 6102 24146
rect 6046 24092 6048 24144
rect 6048 24092 6100 24144
rect 6100 24092 6102 24144
rect 6046 24090 6102 24092
rect 6471 24144 6527 24146
rect 6471 24092 6473 24144
rect 6473 24092 6525 24144
rect 6525 24092 6527 24144
rect 6471 24090 6527 24092
rect 6903 24144 6959 24146
rect 6903 24092 6905 24144
rect 6905 24092 6957 24144
rect 6957 24092 6959 24144
rect 6903 24090 6959 24092
rect 7285 24121 7341 24123
rect 7285 24069 7287 24121
rect 7287 24069 7339 24121
rect 7339 24069 7341 24121
rect 7285 24067 7341 24069
rect 7681 24121 7737 24123
rect 7681 24069 7683 24121
rect 7683 24069 7735 24121
rect 7735 24069 7737 24121
rect 7681 24067 7737 24069
rect 6046 23770 6102 23772
rect 6046 23718 6048 23770
rect 6048 23718 6100 23770
rect 6100 23718 6102 23770
rect 7285 23726 7341 23728
rect 6046 23716 6102 23718
rect 6471 23712 6527 23714
rect 6471 23660 6473 23712
rect 6473 23660 6525 23712
rect 6525 23660 6527 23712
rect 6471 23658 6527 23660
rect 6903 23712 6959 23714
rect 6903 23660 6905 23712
rect 6905 23660 6957 23712
rect 6957 23660 6959 23712
rect 7285 23674 7287 23726
rect 7287 23674 7339 23726
rect 7339 23674 7341 23726
rect 7285 23672 7341 23674
rect 7681 23726 7737 23728
rect 7681 23674 7683 23726
rect 7683 23674 7735 23726
rect 7735 23674 7737 23726
rect 7681 23672 7737 23674
rect 6903 23658 6959 23660
rect 6046 23354 6102 23356
rect 6046 23302 6048 23354
rect 6048 23302 6100 23354
rect 6100 23302 6102 23354
rect 6046 23300 6102 23302
rect 6471 23354 6527 23356
rect 6471 23302 6473 23354
rect 6473 23302 6525 23354
rect 6525 23302 6527 23354
rect 6471 23300 6527 23302
rect 6903 23354 6959 23356
rect 6903 23302 6905 23354
rect 6905 23302 6957 23354
rect 6957 23302 6959 23354
rect 6903 23300 6959 23302
rect 7285 23331 7341 23333
rect 7285 23279 7287 23331
rect 7287 23279 7339 23331
rect 7339 23279 7341 23331
rect 7285 23277 7341 23279
rect 7681 23331 7737 23333
rect 7681 23279 7683 23331
rect 7683 23279 7735 23331
rect 7735 23279 7737 23331
rect 7681 23277 7737 23279
rect 6046 22980 6102 22982
rect 6046 22928 6048 22980
rect 6048 22928 6100 22980
rect 6100 22928 6102 22980
rect 7285 22936 7341 22938
rect 6046 22926 6102 22928
rect 6471 22922 6527 22924
rect 6471 22870 6473 22922
rect 6473 22870 6525 22922
rect 6525 22870 6527 22922
rect 6471 22868 6527 22870
rect 6903 22922 6959 22924
rect 6903 22870 6905 22922
rect 6905 22870 6957 22922
rect 6957 22870 6959 22922
rect 7285 22884 7287 22936
rect 7287 22884 7339 22936
rect 7339 22884 7341 22936
rect 7285 22882 7341 22884
rect 7681 22936 7737 22938
rect 7681 22884 7683 22936
rect 7683 22884 7735 22936
rect 7735 22884 7737 22936
rect 7681 22882 7737 22884
rect 6903 22868 6959 22870
rect 6046 22564 6102 22566
rect 6046 22512 6048 22564
rect 6048 22512 6100 22564
rect 6100 22512 6102 22564
rect 6046 22510 6102 22512
rect 6471 22564 6527 22566
rect 6471 22512 6473 22564
rect 6473 22512 6525 22564
rect 6525 22512 6527 22564
rect 6471 22510 6527 22512
rect 6903 22564 6959 22566
rect 6903 22512 6905 22564
rect 6905 22512 6957 22564
rect 6957 22512 6959 22564
rect 6903 22510 6959 22512
rect 7285 22541 7341 22543
rect 7285 22489 7287 22541
rect 7287 22489 7339 22541
rect 7339 22489 7341 22541
rect 7285 22487 7341 22489
rect 7681 22541 7737 22543
rect 7681 22489 7683 22541
rect 7683 22489 7735 22541
rect 7735 22489 7737 22541
rect 7681 22487 7737 22489
rect 6046 22190 6102 22192
rect 6046 22138 6048 22190
rect 6048 22138 6100 22190
rect 6100 22138 6102 22190
rect 7285 22146 7341 22148
rect 6046 22136 6102 22138
rect 6471 22132 6527 22134
rect 6471 22080 6473 22132
rect 6473 22080 6525 22132
rect 6525 22080 6527 22132
rect 6471 22078 6527 22080
rect 6903 22132 6959 22134
rect 6903 22080 6905 22132
rect 6905 22080 6957 22132
rect 6957 22080 6959 22132
rect 7285 22094 7287 22146
rect 7287 22094 7339 22146
rect 7339 22094 7341 22146
rect 7285 22092 7341 22094
rect 7681 22146 7737 22148
rect 7681 22094 7683 22146
rect 7683 22094 7735 22146
rect 7735 22094 7737 22146
rect 7681 22092 7737 22094
rect 6903 22078 6959 22080
rect 6046 21774 6102 21776
rect 6046 21722 6048 21774
rect 6048 21722 6100 21774
rect 6100 21722 6102 21774
rect 6046 21720 6102 21722
rect 6471 21774 6527 21776
rect 6471 21722 6473 21774
rect 6473 21722 6525 21774
rect 6525 21722 6527 21774
rect 6471 21720 6527 21722
rect 6903 21774 6959 21776
rect 6903 21722 6905 21774
rect 6905 21722 6957 21774
rect 6957 21722 6959 21774
rect 6903 21720 6959 21722
rect 7285 21751 7341 21753
rect 7285 21699 7287 21751
rect 7287 21699 7339 21751
rect 7339 21699 7341 21751
rect 7285 21697 7341 21699
rect 7681 21751 7737 21753
rect 7681 21699 7683 21751
rect 7683 21699 7735 21751
rect 7735 21699 7737 21751
rect 7681 21697 7737 21699
rect 6046 21400 6102 21402
rect 6046 21348 6048 21400
rect 6048 21348 6100 21400
rect 6100 21348 6102 21400
rect 7285 21356 7341 21358
rect 6046 21346 6102 21348
rect 6471 21342 6527 21344
rect 6471 21290 6473 21342
rect 6473 21290 6525 21342
rect 6525 21290 6527 21342
rect 6471 21288 6527 21290
rect 6903 21342 6959 21344
rect 6903 21290 6905 21342
rect 6905 21290 6957 21342
rect 6957 21290 6959 21342
rect 7285 21304 7287 21356
rect 7287 21304 7339 21356
rect 7339 21304 7341 21356
rect 7285 21302 7341 21304
rect 7681 21356 7737 21358
rect 7681 21304 7683 21356
rect 7683 21304 7735 21356
rect 7735 21304 7737 21356
rect 7681 21302 7737 21304
rect 6903 21288 6959 21290
rect 6046 20984 6102 20986
rect 6046 20932 6048 20984
rect 6048 20932 6100 20984
rect 6100 20932 6102 20984
rect 6046 20930 6102 20932
rect 6471 20984 6527 20986
rect 6471 20932 6473 20984
rect 6473 20932 6525 20984
rect 6525 20932 6527 20984
rect 6471 20930 6527 20932
rect 6903 20984 6959 20986
rect 6903 20932 6905 20984
rect 6905 20932 6957 20984
rect 6957 20932 6959 20984
rect 6903 20930 6959 20932
rect 7285 20961 7341 20963
rect 7285 20909 7287 20961
rect 7287 20909 7339 20961
rect 7339 20909 7341 20961
rect 7285 20907 7341 20909
rect 7681 20961 7737 20963
rect 7681 20909 7683 20961
rect 7683 20909 7735 20961
rect 7735 20909 7737 20961
rect 7681 20907 7737 20909
rect 6046 20610 6102 20612
rect 6046 20558 6048 20610
rect 6048 20558 6100 20610
rect 6100 20558 6102 20610
rect 7285 20566 7341 20568
rect 6046 20556 6102 20558
rect 6471 20552 6527 20554
rect 6471 20500 6473 20552
rect 6473 20500 6525 20552
rect 6525 20500 6527 20552
rect 6471 20498 6527 20500
rect 6903 20552 6959 20554
rect 6903 20500 6905 20552
rect 6905 20500 6957 20552
rect 6957 20500 6959 20552
rect 7285 20514 7287 20566
rect 7287 20514 7339 20566
rect 7339 20514 7341 20566
rect 7285 20512 7341 20514
rect 7681 20566 7737 20568
rect 7681 20514 7683 20566
rect 7683 20514 7735 20566
rect 7735 20514 7737 20566
rect 7681 20512 7737 20514
rect 6903 20498 6959 20500
rect 6046 20194 6102 20196
rect 6046 20142 6048 20194
rect 6048 20142 6100 20194
rect 6100 20142 6102 20194
rect 6046 20140 6102 20142
rect 6471 20194 6527 20196
rect 6471 20142 6473 20194
rect 6473 20142 6525 20194
rect 6525 20142 6527 20194
rect 6471 20140 6527 20142
rect 6903 20194 6959 20196
rect 6903 20142 6905 20194
rect 6905 20142 6957 20194
rect 6957 20142 6959 20194
rect 6903 20140 6959 20142
rect 7285 20171 7341 20173
rect 7285 20119 7287 20171
rect 7287 20119 7339 20171
rect 7339 20119 7341 20171
rect 7285 20117 7341 20119
rect 7681 20171 7737 20173
rect 7681 20119 7683 20171
rect 7683 20119 7735 20171
rect 7735 20119 7737 20171
rect 7681 20117 7737 20119
rect 6046 19820 6102 19822
rect 6046 19768 6048 19820
rect 6048 19768 6100 19820
rect 6100 19768 6102 19820
rect 7285 19776 7341 19778
rect 6046 19766 6102 19768
rect 6471 19762 6527 19764
rect 6471 19710 6473 19762
rect 6473 19710 6525 19762
rect 6525 19710 6527 19762
rect 6471 19708 6527 19710
rect 6903 19762 6959 19764
rect 6903 19710 6905 19762
rect 6905 19710 6957 19762
rect 6957 19710 6959 19762
rect 7285 19724 7287 19776
rect 7287 19724 7339 19776
rect 7339 19724 7341 19776
rect 7285 19722 7341 19724
rect 7681 19776 7737 19778
rect 7681 19724 7683 19776
rect 7683 19724 7735 19776
rect 7735 19724 7737 19776
rect 7681 19722 7737 19724
rect 6903 19708 6959 19710
rect 6046 19404 6102 19406
rect 6046 19352 6048 19404
rect 6048 19352 6100 19404
rect 6100 19352 6102 19404
rect 6046 19350 6102 19352
rect 6471 19404 6527 19406
rect 6471 19352 6473 19404
rect 6473 19352 6525 19404
rect 6525 19352 6527 19404
rect 6471 19350 6527 19352
rect 6903 19404 6959 19406
rect 6903 19352 6905 19404
rect 6905 19352 6957 19404
rect 6957 19352 6959 19404
rect 6903 19350 6959 19352
rect 7285 19381 7341 19383
rect 7285 19329 7287 19381
rect 7287 19329 7339 19381
rect 7339 19329 7341 19381
rect 7285 19327 7341 19329
rect 7681 19381 7737 19383
rect 7681 19329 7683 19381
rect 7683 19329 7735 19381
rect 7735 19329 7737 19381
rect 7681 19327 7737 19329
rect 6046 19030 6102 19032
rect 6046 18978 6048 19030
rect 6048 18978 6100 19030
rect 6100 18978 6102 19030
rect 7285 18986 7341 18988
rect 6046 18976 6102 18978
rect 6471 18972 6527 18974
rect 6471 18920 6473 18972
rect 6473 18920 6525 18972
rect 6525 18920 6527 18972
rect 6471 18918 6527 18920
rect 6903 18972 6959 18974
rect 6903 18920 6905 18972
rect 6905 18920 6957 18972
rect 6957 18920 6959 18972
rect 7285 18934 7287 18986
rect 7287 18934 7339 18986
rect 7339 18934 7341 18986
rect 7285 18932 7341 18934
rect 7681 18986 7737 18988
rect 7681 18934 7683 18986
rect 7683 18934 7735 18986
rect 7735 18934 7737 18986
rect 7681 18932 7737 18934
rect 6903 18918 6959 18920
rect 6046 18614 6102 18616
rect 6046 18562 6048 18614
rect 6048 18562 6100 18614
rect 6100 18562 6102 18614
rect 6046 18560 6102 18562
rect 6471 18614 6527 18616
rect 6471 18562 6473 18614
rect 6473 18562 6525 18614
rect 6525 18562 6527 18614
rect 6471 18560 6527 18562
rect 6903 18614 6959 18616
rect 6903 18562 6905 18614
rect 6905 18562 6957 18614
rect 6957 18562 6959 18614
rect 6903 18560 6959 18562
rect 7285 18591 7341 18593
rect 7285 18539 7287 18591
rect 7287 18539 7339 18591
rect 7339 18539 7341 18591
rect 7285 18537 7341 18539
rect 7681 18591 7737 18593
rect 7681 18539 7683 18591
rect 7683 18539 7735 18591
rect 7735 18539 7737 18591
rect 7681 18537 7737 18539
rect 6046 18240 6102 18242
rect 6046 18188 6048 18240
rect 6048 18188 6100 18240
rect 6100 18188 6102 18240
rect 7285 18196 7341 18198
rect 6046 18186 6102 18188
rect 6471 18182 6527 18184
rect 6471 18130 6473 18182
rect 6473 18130 6525 18182
rect 6525 18130 6527 18182
rect 6471 18128 6527 18130
rect 6903 18182 6959 18184
rect 6903 18130 6905 18182
rect 6905 18130 6957 18182
rect 6957 18130 6959 18182
rect 7285 18144 7287 18196
rect 7287 18144 7339 18196
rect 7339 18144 7341 18196
rect 7285 18142 7341 18144
rect 7681 18196 7737 18198
rect 7681 18144 7683 18196
rect 7683 18144 7735 18196
rect 7735 18144 7737 18196
rect 7681 18142 7737 18144
rect 6903 18128 6959 18130
rect 6046 17824 6102 17826
rect 6046 17772 6048 17824
rect 6048 17772 6100 17824
rect 6100 17772 6102 17824
rect 6046 17770 6102 17772
rect 6471 17824 6527 17826
rect 6471 17772 6473 17824
rect 6473 17772 6525 17824
rect 6525 17772 6527 17824
rect 6471 17770 6527 17772
rect 6903 17824 6959 17826
rect 6903 17772 6905 17824
rect 6905 17772 6957 17824
rect 6957 17772 6959 17824
rect 6903 17770 6959 17772
rect 7285 17801 7341 17803
rect 7285 17749 7287 17801
rect 7287 17749 7339 17801
rect 7339 17749 7341 17801
rect 7285 17747 7341 17749
rect 7681 17801 7737 17803
rect 7681 17749 7683 17801
rect 7683 17749 7735 17801
rect 7735 17749 7737 17801
rect 7681 17747 7737 17749
rect 6046 17450 6102 17452
rect 6046 17398 6048 17450
rect 6048 17398 6100 17450
rect 6100 17398 6102 17450
rect 7285 17406 7341 17408
rect 6046 17396 6102 17398
rect 6471 17392 6527 17394
rect 6471 17340 6473 17392
rect 6473 17340 6525 17392
rect 6525 17340 6527 17392
rect 6471 17338 6527 17340
rect 6903 17392 6959 17394
rect 6903 17340 6905 17392
rect 6905 17340 6957 17392
rect 6957 17340 6959 17392
rect 7285 17354 7287 17406
rect 7287 17354 7339 17406
rect 7339 17354 7341 17406
rect 7285 17352 7341 17354
rect 7681 17406 7737 17408
rect 7681 17354 7683 17406
rect 7683 17354 7735 17406
rect 7735 17354 7737 17406
rect 7681 17352 7737 17354
rect 6903 17338 6959 17340
rect 6046 17034 6102 17036
rect 6046 16982 6048 17034
rect 6048 16982 6100 17034
rect 6100 16982 6102 17034
rect 6046 16980 6102 16982
rect 6471 17034 6527 17036
rect 6471 16982 6473 17034
rect 6473 16982 6525 17034
rect 6525 16982 6527 17034
rect 6471 16980 6527 16982
rect 6903 17034 6959 17036
rect 6903 16982 6905 17034
rect 6905 16982 6957 17034
rect 6957 16982 6959 17034
rect 6903 16980 6959 16982
rect 7285 17011 7341 17013
rect 7285 16959 7287 17011
rect 7287 16959 7339 17011
rect 7339 16959 7341 17011
rect 7285 16957 7341 16959
rect 7681 17011 7737 17013
rect 7681 16959 7683 17011
rect 7683 16959 7735 17011
rect 7735 16959 7737 17011
rect 7681 16957 7737 16959
rect 6046 16660 6102 16662
rect 6046 16608 6048 16660
rect 6048 16608 6100 16660
rect 6100 16608 6102 16660
rect 7285 16616 7341 16618
rect 6046 16606 6102 16608
rect 6471 16602 6527 16604
rect 6471 16550 6473 16602
rect 6473 16550 6525 16602
rect 6525 16550 6527 16602
rect 6471 16548 6527 16550
rect 6903 16602 6959 16604
rect 6903 16550 6905 16602
rect 6905 16550 6957 16602
rect 6957 16550 6959 16602
rect 7285 16564 7287 16616
rect 7287 16564 7339 16616
rect 7339 16564 7341 16616
rect 7285 16562 7341 16564
rect 7681 16616 7737 16618
rect 7681 16564 7683 16616
rect 7683 16564 7735 16616
rect 7735 16564 7737 16616
rect 7681 16562 7737 16564
rect 6903 16548 6959 16550
rect 6046 16244 6102 16246
rect 6046 16192 6048 16244
rect 6048 16192 6100 16244
rect 6100 16192 6102 16244
rect 6046 16190 6102 16192
rect 6471 16244 6527 16246
rect 6471 16192 6473 16244
rect 6473 16192 6525 16244
rect 6525 16192 6527 16244
rect 6471 16190 6527 16192
rect 6903 16244 6959 16246
rect 6903 16192 6905 16244
rect 6905 16192 6957 16244
rect 6957 16192 6959 16244
rect 6903 16190 6959 16192
rect 7285 16221 7341 16223
rect 7285 16169 7287 16221
rect 7287 16169 7339 16221
rect 7339 16169 7341 16221
rect 7285 16167 7341 16169
rect 7681 16221 7737 16223
rect 7681 16169 7683 16221
rect 7683 16169 7735 16221
rect 7735 16169 7737 16221
rect 7681 16167 7737 16169
rect 6046 15870 6102 15872
rect 6046 15818 6048 15870
rect 6048 15818 6100 15870
rect 6100 15818 6102 15870
rect 7285 15826 7341 15828
rect 6046 15816 6102 15818
rect 6471 15812 6527 15814
rect 6471 15760 6473 15812
rect 6473 15760 6525 15812
rect 6525 15760 6527 15812
rect 6471 15758 6527 15760
rect 6903 15812 6959 15814
rect 6903 15760 6905 15812
rect 6905 15760 6957 15812
rect 6957 15760 6959 15812
rect 7285 15774 7287 15826
rect 7287 15774 7339 15826
rect 7339 15774 7341 15826
rect 7285 15772 7341 15774
rect 7681 15826 7737 15828
rect 7681 15774 7683 15826
rect 7683 15774 7735 15826
rect 7735 15774 7737 15826
rect 7681 15772 7737 15774
rect 6903 15758 6959 15760
rect 6046 15454 6102 15456
rect 6046 15402 6048 15454
rect 6048 15402 6100 15454
rect 6100 15402 6102 15454
rect 6046 15400 6102 15402
rect 6471 15454 6527 15456
rect 6471 15402 6473 15454
rect 6473 15402 6525 15454
rect 6525 15402 6527 15454
rect 6471 15400 6527 15402
rect 6903 15454 6959 15456
rect 6903 15402 6905 15454
rect 6905 15402 6957 15454
rect 6957 15402 6959 15454
rect 6903 15400 6959 15402
rect 7285 15431 7341 15433
rect 7285 15379 7287 15431
rect 7287 15379 7339 15431
rect 7339 15379 7341 15431
rect 7285 15377 7341 15379
rect 7681 15431 7737 15433
rect 7681 15379 7683 15431
rect 7683 15379 7735 15431
rect 7735 15379 7737 15431
rect 7681 15377 7737 15379
rect 6046 15080 6102 15082
rect 6046 15028 6048 15080
rect 6048 15028 6100 15080
rect 6100 15028 6102 15080
rect 7285 15036 7341 15038
rect 6046 15026 6102 15028
rect 6471 15022 6527 15024
rect 6471 14970 6473 15022
rect 6473 14970 6525 15022
rect 6525 14970 6527 15022
rect 6471 14968 6527 14970
rect 6903 15022 6959 15024
rect 6903 14970 6905 15022
rect 6905 14970 6957 15022
rect 6957 14970 6959 15022
rect 7285 14984 7287 15036
rect 7287 14984 7339 15036
rect 7339 14984 7341 15036
rect 7285 14982 7341 14984
rect 7681 15036 7737 15038
rect 7681 14984 7683 15036
rect 7683 14984 7735 15036
rect 7735 14984 7737 15036
rect 7681 14982 7737 14984
rect 6903 14968 6959 14970
rect 6046 14664 6102 14666
rect 6046 14612 6048 14664
rect 6048 14612 6100 14664
rect 6100 14612 6102 14664
rect 6046 14610 6102 14612
rect 6471 14664 6527 14666
rect 6471 14612 6473 14664
rect 6473 14612 6525 14664
rect 6525 14612 6527 14664
rect 6471 14610 6527 14612
rect 6903 14664 6959 14666
rect 6903 14612 6905 14664
rect 6905 14612 6957 14664
rect 6957 14612 6959 14664
rect 6903 14610 6959 14612
rect 7285 14641 7341 14643
rect 7285 14589 7287 14641
rect 7287 14589 7339 14641
rect 7339 14589 7341 14641
rect 7285 14587 7341 14589
rect 7681 14641 7737 14643
rect 7681 14589 7683 14641
rect 7683 14589 7735 14641
rect 7735 14589 7737 14641
rect 7681 14587 7737 14589
rect 6046 14290 6102 14292
rect 6046 14238 6048 14290
rect 6048 14238 6100 14290
rect 6100 14238 6102 14290
rect 7285 14246 7341 14248
rect 6046 14236 6102 14238
rect 6471 14232 6527 14234
rect 6471 14180 6473 14232
rect 6473 14180 6525 14232
rect 6525 14180 6527 14232
rect 6471 14178 6527 14180
rect 6903 14232 6959 14234
rect 6903 14180 6905 14232
rect 6905 14180 6957 14232
rect 6957 14180 6959 14232
rect 7285 14194 7287 14246
rect 7287 14194 7339 14246
rect 7339 14194 7341 14246
rect 7285 14192 7341 14194
rect 7681 14246 7737 14248
rect 7681 14194 7683 14246
rect 7683 14194 7735 14246
rect 7735 14194 7737 14246
rect 7681 14192 7737 14194
rect 6903 14178 6959 14180
rect 6046 13874 6102 13876
rect 6046 13822 6048 13874
rect 6048 13822 6100 13874
rect 6100 13822 6102 13874
rect 6046 13820 6102 13822
rect 6471 13874 6527 13876
rect 6471 13822 6473 13874
rect 6473 13822 6525 13874
rect 6525 13822 6527 13874
rect 6471 13820 6527 13822
rect 6903 13874 6959 13876
rect 6903 13822 6905 13874
rect 6905 13822 6957 13874
rect 6957 13822 6959 13874
rect 6903 13820 6959 13822
rect 7285 13851 7341 13853
rect 7285 13799 7287 13851
rect 7287 13799 7339 13851
rect 7339 13799 7341 13851
rect 7285 13797 7341 13799
rect 7681 13851 7737 13853
rect 7681 13799 7683 13851
rect 7683 13799 7735 13851
rect 7735 13799 7737 13851
rect 7681 13797 7737 13799
rect 6046 13500 6102 13502
rect 6046 13448 6048 13500
rect 6048 13448 6100 13500
rect 6100 13448 6102 13500
rect 7285 13456 7341 13458
rect 6046 13446 6102 13448
rect 6471 13442 6527 13444
rect 6471 13390 6473 13442
rect 6473 13390 6525 13442
rect 6525 13390 6527 13442
rect 6471 13388 6527 13390
rect 6903 13442 6959 13444
rect 6903 13390 6905 13442
rect 6905 13390 6957 13442
rect 6957 13390 6959 13442
rect 7285 13404 7287 13456
rect 7287 13404 7339 13456
rect 7339 13404 7341 13456
rect 7285 13402 7341 13404
rect 7681 13456 7737 13458
rect 7681 13404 7683 13456
rect 7683 13404 7735 13456
rect 7735 13404 7737 13456
rect 7681 13402 7737 13404
rect 6903 13388 6959 13390
rect 6046 13084 6102 13086
rect 6046 13032 6048 13084
rect 6048 13032 6100 13084
rect 6100 13032 6102 13084
rect 6046 13030 6102 13032
rect 6471 13084 6527 13086
rect 6471 13032 6473 13084
rect 6473 13032 6525 13084
rect 6525 13032 6527 13084
rect 6471 13030 6527 13032
rect 6903 13084 6959 13086
rect 6903 13032 6905 13084
rect 6905 13032 6957 13084
rect 6957 13032 6959 13084
rect 6903 13030 6959 13032
rect 7285 13061 7341 13063
rect 7285 13009 7287 13061
rect 7287 13009 7339 13061
rect 7339 13009 7341 13061
rect 7285 13007 7341 13009
rect 7681 13061 7737 13063
rect 7681 13009 7683 13061
rect 7683 13009 7735 13061
rect 7735 13009 7737 13061
rect 7681 13007 7737 13009
rect 6046 12710 6102 12712
rect 6046 12658 6048 12710
rect 6048 12658 6100 12710
rect 6100 12658 6102 12710
rect 7285 12666 7341 12668
rect 6046 12656 6102 12658
rect 6471 12652 6527 12654
rect 6471 12600 6473 12652
rect 6473 12600 6525 12652
rect 6525 12600 6527 12652
rect 6471 12598 6527 12600
rect 6903 12652 6959 12654
rect 6903 12600 6905 12652
rect 6905 12600 6957 12652
rect 6957 12600 6959 12652
rect 7285 12614 7287 12666
rect 7287 12614 7339 12666
rect 7339 12614 7341 12666
rect 7285 12612 7341 12614
rect 7681 12666 7737 12668
rect 7681 12614 7683 12666
rect 7683 12614 7735 12666
rect 7735 12614 7737 12666
rect 7681 12612 7737 12614
rect 6903 12598 6959 12600
rect 6046 12294 6102 12296
rect 6046 12242 6048 12294
rect 6048 12242 6100 12294
rect 6100 12242 6102 12294
rect 6046 12240 6102 12242
rect 6471 12294 6527 12296
rect 6471 12242 6473 12294
rect 6473 12242 6525 12294
rect 6525 12242 6527 12294
rect 6471 12240 6527 12242
rect 6903 12294 6959 12296
rect 6903 12242 6905 12294
rect 6905 12242 6957 12294
rect 6957 12242 6959 12294
rect 6903 12240 6959 12242
rect 7285 12271 7341 12273
rect 7285 12219 7287 12271
rect 7287 12219 7339 12271
rect 7339 12219 7341 12271
rect 7285 12217 7341 12219
rect 7681 12271 7737 12273
rect 7681 12219 7683 12271
rect 7683 12219 7735 12271
rect 7735 12219 7737 12271
rect 7681 12217 7737 12219
rect 6046 11920 6102 11922
rect 6046 11868 6048 11920
rect 6048 11868 6100 11920
rect 6100 11868 6102 11920
rect 7285 11876 7341 11878
rect 6046 11866 6102 11868
rect 6471 11862 6527 11864
rect 6471 11810 6473 11862
rect 6473 11810 6525 11862
rect 6525 11810 6527 11862
rect 6471 11808 6527 11810
rect 6903 11862 6959 11864
rect 6903 11810 6905 11862
rect 6905 11810 6957 11862
rect 6957 11810 6959 11862
rect 7285 11824 7287 11876
rect 7287 11824 7339 11876
rect 7339 11824 7341 11876
rect 7285 11822 7341 11824
rect 7681 11876 7737 11878
rect 7681 11824 7683 11876
rect 7683 11824 7735 11876
rect 7735 11824 7737 11876
rect 7681 11822 7737 11824
rect 6903 11808 6959 11810
rect 6046 11504 6102 11506
rect 6046 11452 6048 11504
rect 6048 11452 6100 11504
rect 6100 11452 6102 11504
rect 6046 11450 6102 11452
rect 6471 11504 6527 11506
rect 6471 11452 6473 11504
rect 6473 11452 6525 11504
rect 6525 11452 6527 11504
rect 6471 11450 6527 11452
rect 6903 11504 6959 11506
rect 6903 11452 6905 11504
rect 6905 11452 6957 11504
rect 6957 11452 6959 11504
rect 6903 11450 6959 11452
rect 7285 11481 7341 11483
rect 7285 11429 7287 11481
rect 7287 11429 7339 11481
rect 7339 11429 7341 11481
rect 7285 11427 7341 11429
rect 7681 11481 7737 11483
rect 7681 11429 7683 11481
rect 7683 11429 7735 11481
rect 7735 11429 7737 11481
rect 7681 11427 7737 11429
rect 6046 11130 6102 11132
rect 6046 11078 6048 11130
rect 6048 11078 6100 11130
rect 6100 11078 6102 11130
rect 7285 11086 7341 11088
rect 6046 11076 6102 11078
rect 6471 11072 6527 11074
rect 6471 11020 6473 11072
rect 6473 11020 6525 11072
rect 6525 11020 6527 11072
rect 6471 11018 6527 11020
rect 6903 11072 6959 11074
rect 6903 11020 6905 11072
rect 6905 11020 6957 11072
rect 6957 11020 6959 11072
rect 7285 11034 7287 11086
rect 7287 11034 7339 11086
rect 7339 11034 7341 11086
rect 7285 11032 7341 11034
rect 7681 11086 7737 11088
rect 7681 11034 7683 11086
rect 7683 11034 7735 11086
rect 7735 11034 7737 11086
rect 7681 11032 7737 11034
rect 6903 11018 6959 11020
rect 6046 10714 6102 10716
rect 6046 10662 6048 10714
rect 6048 10662 6100 10714
rect 6100 10662 6102 10714
rect 6046 10660 6102 10662
rect 6471 10714 6527 10716
rect 6471 10662 6473 10714
rect 6473 10662 6525 10714
rect 6525 10662 6527 10714
rect 6471 10660 6527 10662
rect 6903 10714 6959 10716
rect 6903 10662 6905 10714
rect 6905 10662 6957 10714
rect 6957 10662 6959 10714
rect 6903 10660 6959 10662
rect 7285 10691 7341 10693
rect 7285 10639 7287 10691
rect 7287 10639 7339 10691
rect 7339 10639 7341 10691
rect 7285 10637 7341 10639
rect 7681 10691 7737 10693
rect 7681 10639 7683 10691
rect 7683 10639 7735 10691
rect 7735 10639 7737 10691
rect 7681 10637 7737 10639
rect 6046 10340 6102 10342
rect 6046 10288 6048 10340
rect 6048 10288 6100 10340
rect 6100 10288 6102 10340
rect 7285 10296 7341 10298
rect 6046 10286 6102 10288
rect 6471 10282 6527 10284
rect 6471 10230 6473 10282
rect 6473 10230 6525 10282
rect 6525 10230 6527 10282
rect 6471 10228 6527 10230
rect 6903 10282 6959 10284
rect 6903 10230 6905 10282
rect 6905 10230 6957 10282
rect 6957 10230 6959 10282
rect 7285 10244 7287 10296
rect 7287 10244 7339 10296
rect 7339 10244 7341 10296
rect 7285 10242 7341 10244
rect 7681 10296 7737 10298
rect 7681 10244 7683 10296
rect 7683 10244 7735 10296
rect 7735 10244 7737 10296
rect 7681 10242 7737 10244
rect 6903 10228 6959 10230
rect 6046 9924 6102 9926
rect 6046 9872 6048 9924
rect 6048 9872 6100 9924
rect 6100 9872 6102 9924
rect 6046 9870 6102 9872
rect 6471 9924 6527 9926
rect 6471 9872 6473 9924
rect 6473 9872 6525 9924
rect 6525 9872 6527 9924
rect 6471 9870 6527 9872
rect 6903 9924 6959 9926
rect 6903 9872 6905 9924
rect 6905 9872 6957 9924
rect 6957 9872 6959 9924
rect 6903 9870 6959 9872
rect 7285 9901 7341 9903
rect 7285 9849 7287 9901
rect 7287 9849 7339 9901
rect 7339 9849 7341 9901
rect 7285 9847 7341 9849
rect 7681 9901 7737 9903
rect 7681 9849 7683 9901
rect 7683 9849 7735 9901
rect 7735 9849 7737 9901
rect 7681 9847 7737 9849
rect 6046 9550 6102 9552
rect 6046 9498 6048 9550
rect 6048 9498 6100 9550
rect 6100 9498 6102 9550
rect 7285 9506 7341 9508
rect 6046 9496 6102 9498
rect 6471 9492 6527 9494
rect 6471 9440 6473 9492
rect 6473 9440 6525 9492
rect 6525 9440 6527 9492
rect 6471 9438 6527 9440
rect 6903 9492 6959 9494
rect 6903 9440 6905 9492
rect 6905 9440 6957 9492
rect 6957 9440 6959 9492
rect 7285 9454 7287 9506
rect 7287 9454 7339 9506
rect 7339 9454 7341 9506
rect 7285 9452 7341 9454
rect 7681 9506 7737 9508
rect 7681 9454 7683 9506
rect 7683 9454 7735 9506
rect 7735 9454 7737 9506
rect 7681 9452 7737 9454
rect 6903 9438 6959 9440
rect 6046 9134 6102 9136
rect 6046 9082 6048 9134
rect 6048 9082 6100 9134
rect 6100 9082 6102 9134
rect 6046 9080 6102 9082
rect 6471 9134 6527 9136
rect 6471 9082 6473 9134
rect 6473 9082 6525 9134
rect 6525 9082 6527 9134
rect 6471 9080 6527 9082
rect 6903 9134 6959 9136
rect 6903 9082 6905 9134
rect 6905 9082 6957 9134
rect 6957 9082 6959 9134
rect 6903 9080 6959 9082
rect 7285 9111 7341 9113
rect 7285 9059 7287 9111
rect 7287 9059 7339 9111
rect 7339 9059 7341 9111
rect 7285 9057 7341 9059
rect 7681 9111 7737 9113
rect 7681 9059 7683 9111
rect 7683 9059 7735 9111
rect 7735 9059 7737 9111
rect 7681 9057 7737 9059
rect 6046 8760 6102 8762
rect 6046 8708 6048 8760
rect 6048 8708 6100 8760
rect 6100 8708 6102 8760
rect 7285 8716 7341 8718
rect 6046 8706 6102 8708
rect 6471 8702 6527 8704
rect 6471 8650 6473 8702
rect 6473 8650 6525 8702
rect 6525 8650 6527 8702
rect 6471 8648 6527 8650
rect 6903 8702 6959 8704
rect 6903 8650 6905 8702
rect 6905 8650 6957 8702
rect 6957 8650 6959 8702
rect 7285 8664 7287 8716
rect 7287 8664 7339 8716
rect 7339 8664 7341 8716
rect 7285 8662 7341 8664
rect 7681 8716 7737 8718
rect 7681 8664 7683 8716
rect 7683 8664 7735 8716
rect 7735 8664 7737 8716
rect 7681 8662 7737 8664
rect 6903 8648 6959 8650
rect 6046 8344 6102 8346
rect 6046 8292 6048 8344
rect 6048 8292 6100 8344
rect 6100 8292 6102 8344
rect 6046 8290 6102 8292
rect 6471 8344 6527 8346
rect 6471 8292 6473 8344
rect 6473 8292 6525 8344
rect 6525 8292 6527 8344
rect 6471 8290 6527 8292
rect 6903 8344 6959 8346
rect 6903 8292 6905 8344
rect 6905 8292 6957 8344
rect 6957 8292 6959 8344
rect 6903 8290 6959 8292
rect 7285 8321 7341 8323
rect 7285 8269 7287 8321
rect 7287 8269 7339 8321
rect 7339 8269 7341 8321
rect 7285 8267 7341 8269
rect 7681 8321 7737 8323
rect 7681 8269 7683 8321
rect 7683 8269 7735 8321
rect 7735 8269 7737 8321
rect 7681 8267 7737 8269
rect 6046 7970 6102 7972
rect 6046 7918 6048 7970
rect 6048 7918 6100 7970
rect 6100 7918 6102 7970
rect 7285 7926 7341 7928
rect 6046 7916 6102 7918
rect 6471 7912 6527 7914
rect 6471 7860 6473 7912
rect 6473 7860 6525 7912
rect 6525 7860 6527 7912
rect 6471 7858 6527 7860
rect 6903 7912 6959 7914
rect 6903 7860 6905 7912
rect 6905 7860 6957 7912
rect 6957 7860 6959 7912
rect 7285 7874 7287 7926
rect 7287 7874 7339 7926
rect 7339 7874 7341 7926
rect 7285 7872 7341 7874
rect 7681 7926 7737 7928
rect 7681 7874 7683 7926
rect 7683 7874 7735 7926
rect 7735 7874 7737 7926
rect 7681 7872 7737 7874
rect 6903 7858 6959 7860
rect 6046 7554 6102 7556
rect 6046 7502 6048 7554
rect 6048 7502 6100 7554
rect 6100 7502 6102 7554
rect 6046 7500 6102 7502
rect 6471 7554 6527 7556
rect 6471 7502 6473 7554
rect 6473 7502 6525 7554
rect 6525 7502 6527 7554
rect 6471 7500 6527 7502
rect 6903 7554 6959 7556
rect 6903 7502 6905 7554
rect 6905 7502 6957 7554
rect 6957 7502 6959 7554
rect 6903 7500 6959 7502
rect 7285 7531 7341 7533
rect 7285 7479 7287 7531
rect 7287 7479 7339 7531
rect 7339 7479 7341 7531
rect 7285 7477 7341 7479
rect 7681 7531 7737 7533
rect 7681 7479 7683 7531
rect 7683 7479 7735 7531
rect 7735 7479 7737 7531
rect 7681 7477 7737 7479
rect 6046 7180 6102 7182
rect 6046 7128 6048 7180
rect 6048 7128 6100 7180
rect 6100 7128 6102 7180
rect 7285 7136 7341 7138
rect 6046 7126 6102 7128
rect 6471 7122 6527 7124
rect 6471 7070 6473 7122
rect 6473 7070 6525 7122
rect 6525 7070 6527 7122
rect 6471 7068 6527 7070
rect 6903 7122 6959 7124
rect 6903 7070 6905 7122
rect 6905 7070 6957 7122
rect 6957 7070 6959 7122
rect 7285 7084 7287 7136
rect 7287 7084 7339 7136
rect 7339 7084 7341 7136
rect 7285 7082 7341 7084
rect 7681 7136 7737 7138
rect 7681 7084 7683 7136
rect 7683 7084 7735 7136
rect 7735 7084 7737 7136
rect 7681 7082 7737 7084
rect 6903 7068 6959 7070
rect 6046 6764 6102 6766
rect 6046 6712 6048 6764
rect 6048 6712 6100 6764
rect 6100 6712 6102 6764
rect 6046 6710 6102 6712
rect 6471 6764 6527 6766
rect 6471 6712 6473 6764
rect 6473 6712 6525 6764
rect 6525 6712 6527 6764
rect 6471 6710 6527 6712
rect 6903 6764 6959 6766
rect 6903 6712 6905 6764
rect 6905 6712 6957 6764
rect 6957 6712 6959 6764
rect 6903 6710 6959 6712
rect 7285 6741 7341 6743
rect 7285 6689 7287 6741
rect 7287 6689 7339 6741
rect 7339 6689 7341 6741
rect 7285 6687 7341 6689
rect 7681 6741 7737 6743
rect 7681 6689 7683 6741
rect 7683 6689 7735 6741
rect 7735 6689 7737 6741
rect 7681 6687 7737 6689
rect 6046 6390 6102 6392
rect 6046 6338 6048 6390
rect 6048 6338 6100 6390
rect 6100 6338 6102 6390
rect 7285 6346 7341 6348
rect 6046 6336 6102 6338
rect 6471 6332 6527 6334
rect 6471 6280 6473 6332
rect 6473 6280 6525 6332
rect 6525 6280 6527 6332
rect 6471 6278 6527 6280
rect 6903 6332 6959 6334
rect 6903 6280 6905 6332
rect 6905 6280 6957 6332
rect 6957 6280 6959 6332
rect 7285 6294 7287 6346
rect 7287 6294 7339 6346
rect 7339 6294 7341 6346
rect 7285 6292 7341 6294
rect 7681 6346 7737 6348
rect 7681 6294 7683 6346
rect 7683 6294 7735 6346
rect 7735 6294 7737 6346
rect 7681 6292 7737 6294
rect 6903 6278 6959 6280
rect 6046 5974 6102 5976
rect 6046 5922 6048 5974
rect 6048 5922 6100 5974
rect 6100 5922 6102 5974
rect 6046 5920 6102 5922
rect 6471 5974 6527 5976
rect 6471 5922 6473 5974
rect 6473 5922 6525 5974
rect 6525 5922 6527 5974
rect 6471 5920 6527 5922
rect 6903 5974 6959 5976
rect 6903 5922 6905 5974
rect 6905 5922 6957 5974
rect 6957 5922 6959 5974
rect 6903 5920 6959 5922
rect 7285 5951 7341 5953
rect 7285 5899 7287 5951
rect 7287 5899 7339 5951
rect 7339 5899 7341 5951
rect 7285 5897 7341 5899
rect 7681 5951 7737 5953
rect 7681 5899 7683 5951
rect 7683 5899 7735 5951
rect 7735 5899 7737 5951
rect 7681 5897 7737 5899
rect 6046 5600 6102 5602
rect 6046 5548 6048 5600
rect 6048 5548 6100 5600
rect 6100 5548 6102 5600
rect 7285 5556 7341 5558
rect 6046 5546 6102 5548
rect 6471 5542 6527 5544
rect 6471 5490 6473 5542
rect 6473 5490 6525 5542
rect 6525 5490 6527 5542
rect 6471 5488 6527 5490
rect 6903 5542 6959 5544
rect 6903 5490 6905 5542
rect 6905 5490 6957 5542
rect 6957 5490 6959 5542
rect 7285 5504 7287 5556
rect 7287 5504 7339 5556
rect 7339 5504 7341 5556
rect 7285 5502 7341 5504
rect 7681 5556 7737 5558
rect 7681 5504 7683 5556
rect 7683 5504 7735 5556
rect 7735 5504 7737 5556
rect 7681 5502 7737 5504
rect 6903 5488 6959 5490
rect 6046 5184 6102 5186
rect 6046 5132 6048 5184
rect 6048 5132 6100 5184
rect 6100 5132 6102 5184
rect 6046 5130 6102 5132
rect 6471 5184 6527 5186
rect 6471 5132 6473 5184
rect 6473 5132 6525 5184
rect 6525 5132 6527 5184
rect 6471 5130 6527 5132
rect 6903 5184 6959 5186
rect 6903 5132 6905 5184
rect 6905 5132 6957 5184
rect 6957 5132 6959 5184
rect 6903 5130 6959 5132
rect 7285 5161 7341 5163
rect 7285 5109 7287 5161
rect 7287 5109 7339 5161
rect 7339 5109 7341 5161
rect 7285 5107 7341 5109
rect 7681 5161 7737 5163
rect 7681 5109 7683 5161
rect 7683 5109 7735 5161
rect 7735 5109 7737 5161
rect 7681 5107 7737 5109
rect 6046 4810 6102 4812
rect 6046 4758 6048 4810
rect 6048 4758 6100 4810
rect 6100 4758 6102 4810
rect 7285 4766 7341 4768
rect 6046 4756 6102 4758
rect 6471 4752 6527 4754
rect 6471 4700 6473 4752
rect 6473 4700 6525 4752
rect 6525 4700 6527 4752
rect 6471 4698 6527 4700
rect 6903 4752 6959 4754
rect 6903 4700 6905 4752
rect 6905 4700 6957 4752
rect 6957 4700 6959 4752
rect 7285 4714 7287 4766
rect 7287 4714 7339 4766
rect 7339 4714 7341 4766
rect 7285 4712 7341 4714
rect 7681 4766 7737 4768
rect 7681 4714 7683 4766
rect 7683 4714 7735 4766
rect 7735 4714 7737 4766
rect 7681 4712 7737 4714
rect 6903 4698 6959 4700
rect 6046 4394 6102 4396
rect 6046 4342 6048 4394
rect 6048 4342 6100 4394
rect 6100 4342 6102 4394
rect 6046 4340 6102 4342
rect 6471 4394 6527 4396
rect 6471 4342 6473 4394
rect 6473 4342 6525 4394
rect 6525 4342 6527 4394
rect 6471 4340 6527 4342
rect 6903 4394 6959 4396
rect 6903 4342 6905 4394
rect 6905 4342 6957 4394
rect 6957 4342 6959 4394
rect 6903 4340 6959 4342
rect 7285 4371 7341 4373
rect 7285 4319 7287 4371
rect 7287 4319 7339 4371
rect 7339 4319 7341 4371
rect 7285 4317 7341 4319
rect 7681 4371 7737 4373
rect 7681 4319 7683 4371
rect 7683 4319 7735 4371
rect 7735 4319 7737 4371
rect 7681 4317 7737 4319
rect 6046 4020 6102 4022
rect 6046 3968 6048 4020
rect 6048 3968 6100 4020
rect 6100 3968 6102 4020
rect 7285 3976 7341 3978
rect 6046 3966 6102 3968
rect 6471 3962 6527 3964
rect 6471 3910 6473 3962
rect 6473 3910 6525 3962
rect 6525 3910 6527 3962
rect 6471 3908 6527 3910
rect 6903 3962 6959 3964
rect 6903 3910 6905 3962
rect 6905 3910 6957 3962
rect 6957 3910 6959 3962
rect 7285 3924 7287 3976
rect 7287 3924 7339 3976
rect 7339 3924 7341 3976
rect 7285 3922 7341 3924
rect 7681 3976 7737 3978
rect 7681 3924 7683 3976
rect 7683 3924 7735 3976
rect 7735 3924 7737 3976
rect 7681 3922 7737 3924
rect 6903 3908 6959 3910
rect 6046 3604 6102 3606
rect 6046 3552 6048 3604
rect 6048 3552 6100 3604
rect 6100 3552 6102 3604
rect 6046 3550 6102 3552
rect 6471 3604 6527 3606
rect 6471 3552 6473 3604
rect 6473 3552 6525 3604
rect 6525 3552 6527 3604
rect 6471 3550 6527 3552
rect 6903 3604 6959 3606
rect 6903 3552 6905 3604
rect 6905 3552 6957 3604
rect 6957 3552 6959 3604
rect 6903 3550 6959 3552
rect 7285 3581 7341 3583
rect 7285 3529 7287 3581
rect 7287 3529 7339 3581
rect 7339 3529 7341 3581
rect 7285 3527 7341 3529
rect 7681 3581 7737 3583
rect 7681 3529 7683 3581
rect 7683 3529 7735 3581
rect 7735 3529 7737 3581
rect 7681 3527 7737 3529
rect 6046 3230 6102 3232
rect 6046 3178 6048 3230
rect 6048 3178 6100 3230
rect 6100 3178 6102 3230
rect 7285 3186 7341 3188
rect 6046 3176 6102 3178
rect 6471 3172 6527 3174
rect 6471 3120 6473 3172
rect 6473 3120 6525 3172
rect 6525 3120 6527 3172
rect 6471 3118 6527 3120
rect 6903 3172 6959 3174
rect 6903 3120 6905 3172
rect 6905 3120 6957 3172
rect 6957 3120 6959 3172
rect 7285 3134 7287 3186
rect 7287 3134 7339 3186
rect 7339 3134 7341 3186
rect 7285 3132 7341 3134
rect 7681 3186 7737 3188
rect 7681 3134 7683 3186
rect 7683 3134 7735 3186
rect 7735 3134 7737 3186
rect 7681 3132 7737 3134
rect 6903 3118 6959 3120
rect 6046 2814 6102 2816
rect 6046 2762 6048 2814
rect 6048 2762 6100 2814
rect 6100 2762 6102 2814
rect 6046 2760 6102 2762
rect 6471 2814 6527 2816
rect 6471 2762 6473 2814
rect 6473 2762 6525 2814
rect 6525 2762 6527 2814
rect 6471 2760 6527 2762
rect 6903 2814 6959 2816
rect 6903 2762 6905 2814
rect 6905 2762 6957 2814
rect 6957 2762 6959 2814
rect 6903 2760 6959 2762
rect 7285 2791 7341 2793
rect 7285 2739 7287 2791
rect 7287 2739 7339 2791
rect 7339 2739 7341 2791
rect 7285 2737 7341 2739
rect 7681 2791 7737 2793
rect 7681 2739 7683 2791
rect 7683 2739 7735 2791
rect 7735 2739 7737 2791
rect 7681 2737 7737 2739
rect 6046 2440 6102 2442
rect 6046 2388 6048 2440
rect 6048 2388 6100 2440
rect 6100 2388 6102 2440
rect 7285 2396 7341 2398
rect 6046 2386 6102 2388
rect 6471 2382 6527 2384
rect 6471 2330 6473 2382
rect 6473 2330 6525 2382
rect 6525 2330 6527 2382
rect 6471 2328 6527 2330
rect 6903 2382 6959 2384
rect 6903 2330 6905 2382
rect 6905 2330 6957 2382
rect 6957 2330 6959 2382
rect 7285 2344 7287 2396
rect 7287 2344 7339 2396
rect 7339 2344 7341 2396
rect 7285 2342 7341 2344
rect 7681 2396 7737 2398
rect 7681 2344 7683 2396
rect 7683 2344 7735 2396
rect 7735 2344 7737 2396
rect 7681 2342 7737 2344
rect 6903 2328 6959 2330
rect 6046 2024 6102 2026
rect 6046 1972 6048 2024
rect 6048 1972 6100 2024
rect 6100 1972 6102 2024
rect 6046 1970 6102 1972
rect 6471 2024 6527 2026
rect 6471 1972 6473 2024
rect 6473 1972 6525 2024
rect 6525 1972 6527 2024
rect 6471 1970 6527 1972
rect 6903 2024 6959 2026
rect 6903 1972 6905 2024
rect 6905 1972 6957 2024
rect 6957 1972 6959 2024
rect 6903 1970 6959 1972
rect 7285 2001 7341 2003
rect 7285 1949 7287 2001
rect 7287 1949 7339 2001
rect 7339 1949 7341 2001
rect 7285 1947 7341 1949
rect 7681 2001 7737 2003
rect 7681 1949 7683 2001
rect 7683 1949 7735 2001
rect 7735 1949 7737 2001
rect 7681 1947 7737 1949
rect 6046 1650 6102 1652
rect 6046 1598 6048 1650
rect 6048 1598 6100 1650
rect 6100 1598 6102 1650
rect 7285 1606 7341 1608
rect 6046 1596 6102 1598
rect 6471 1592 6527 1594
rect 6471 1540 6473 1592
rect 6473 1540 6525 1592
rect 6525 1540 6527 1592
rect 6471 1538 6527 1540
rect 6903 1592 6959 1594
rect 6903 1540 6905 1592
rect 6905 1540 6957 1592
rect 6957 1540 6959 1592
rect 7285 1554 7287 1606
rect 7287 1554 7339 1606
rect 7339 1554 7341 1606
rect 7285 1552 7341 1554
rect 7681 1606 7737 1608
rect 7681 1554 7683 1606
rect 7683 1554 7735 1606
rect 7735 1554 7737 1606
rect 7681 1552 7737 1554
rect 6903 1538 6959 1540
rect 6046 1234 6102 1236
rect 6046 1182 6048 1234
rect 6048 1182 6100 1234
rect 6100 1182 6102 1234
rect 6046 1180 6102 1182
rect 6471 1234 6527 1236
rect 6471 1182 6473 1234
rect 6473 1182 6525 1234
rect 6525 1182 6527 1234
rect 6471 1180 6527 1182
rect 6903 1234 6959 1236
rect 6903 1182 6905 1234
rect 6905 1182 6957 1234
rect 6957 1182 6959 1234
rect 6903 1180 6959 1182
rect 7285 1211 7341 1213
rect 7285 1159 7287 1211
rect 7287 1159 7339 1211
rect 7339 1159 7341 1211
rect 7285 1157 7341 1159
rect 7681 1211 7737 1213
rect 7681 1159 7683 1211
rect 7683 1159 7735 1211
rect 7735 1159 7737 1211
rect 7681 1157 7737 1159
rect 6046 860 6102 862
rect 6046 808 6048 860
rect 6048 808 6100 860
rect 6100 808 6102 860
rect 7285 816 7341 818
rect 6046 806 6102 808
rect 6471 802 6527 804
rect 6471 750 6473 802
rect 6473 750 6525 802
rect 6525 750 6527 802
rect 6471 748 6527 750
rect 6903 802 6959 804
rect 6903 750 6905 802
rect 6905 750 6957 802
rect 6957 750 6959 802
rect 7285 764 7287 816
rect 7287 764 7339 816
rect 7339 764 7341 816
rect 7285 762 7341 764
rect 7681 816 7737 818
rect 7681 764 7683 816
rect 7683 764 7735 816
rect 7735 764 7737 816
rect 7681 762 7737 764
rect 6903 748 6959 750
rect 6046 444 6102 446
rect 6046 392 6048 444
rect 6048 392 6100 444
rect 6100 392 6102 444
rect 6046 390 6102 392
rect 6471 444 6527 446
rect 6471 392 6473 444
rect 6473 392 6525 444
rect 6525 392 6527 444
rect 6471 390 6527 392
rect 6903 444 6959 446
rect 6903 392 6905 444
rect 6905 392 6957 444
rect 6957 392 6959 444
rect 6903 390 6959 392
rect 7285 421 7341 423
rect 7285 369 7287 421
rect 7287 369 7339 421
rect 7339 369 7341 421
rect 7285 367 7341 369
rect 7681 421 7737 423
rect 7681 369 7683 421
rect 7683 369 7735 421
rect 7735 369 7737 421
rect 7681 367 7737 369
<< metal3 >>
rect 6025 50216 6123 50237
rect 6025 50160 6046 50216
rect 6102 50160 6123 50216
rect 6025 50139 6123 50160
rect 6450 50216 6548 50237
rect 6450 50160 6471 50216
rect 6527 50160 6548 50216
rect 6450 50139 6548 50160
rect 6882 50216 6980 50237
rect 6882 50160 6903 50216
rect 6959 50160 6980 50216
rect 6882 50139 6980 50160
rect 7264 50193 7362 50214
rect 7264 50137 7285 50193
rect 7341 50137 7362 50193
rect 7264 50116 7362 50137
rect 7660 50193 7758 50214
rect 7660 50137 7681 50193
rect 7737 50137 7758 50193
rect 7660 50116 7758 50137
rect 6025 49842 6123 49863
rect 6025 49786 6046 49842
rect 6102 49786 6123 49842
rect 6025 49765 6123 49786
rect 6450 49784 6548 49805
rect 6450 49728 6471 49784
rect 6527 49728 6548 49784
rect 6450 49707 6548 49728
rect 6882 49784 6980 49805
rect 6882 49728 6903 49784
rect 6959 49728 6980 49784
rect 6882 49707 6980 49728
rect 7264 49798 7362 49819
rect 7264 49742 7285 49798
rect 7341 49742 7362 49798
rect 7264 49721 7362 49742
rect 7660 49798 7758 49819
rect 7660 49742 7681 49798
rect 7737 49742 7758 49798
rect 7660 49721 7758 49742
rect 6025 49426 6123 49447
rect 6025 49370 6046 49426
rect 6102 49370 6123 49426
rect 6025 49349 6123 49370
rect 6450 49426 6548 49447
rect 6450 49370 6471 49426
rect 6527 49370 6548 49426
rect 6450 49349 6548 49370
rect 6882 49426 6980 49447
rect 6882 49370 6903 49426
rect 6959 49370 6980 49426
rect 6882 49349 6980 49370
rect 7264 49403 7362 49424
rect 7264 49347 7285 49403
rect 7341 49347 7362 49403
rect 7264 49326 7362 49347
rect 7660 49403 7758 49424
rect 7660 49347 7681 49403
rect 7737 49347 7758 49403
rect 7660 49326 7758 49347
rect 6025 49052 6123 49073
rect 6025 48996 6046 49052
rect 6102 48996 6123 49052
rect 6025 48975 6123 48996
rect 6450 48994 6548 49015
rect 6450 48938 6471 48994
rect 6527 48938 6548 48994
rect 6450 48917 6548 48938
rect 6882 48994 6980 49015
rect 6882 48938 6903 48994
rect 6959 48938 6980 48994
rect 6882 48917 6980 48938
rect 7264 49008 7362 49029
rect 7264 48952 7285 49008
rect 7341 48952 7362 49008
rect 7264 48931 7362 48952
rect 7660 49008 7758 49029
rect 7660 48952 7681 49008
rect 7737 48952 7758 49008
rect 7660 48931 7758 48952
rect 6025 48636 6123 48657
rect 6025 48580 6046 48636
rect 6102 48580 6123 48636
rect 6025 48559 6123 48580
rect 6450 48636 6548 48657
rect 6450 48580 6471 48636
rect 6527 48580 6548 48636
rect 6450 48559 6548 48580
rect 6882 48636 6980 48657
rect 6882 48580 6903 48636
rect 6959 48580 6980 48636
rect 6882 48559 6980 48580
rect 7264 48613 7362 48634
rect 7264 48557 7285 48613
rect 7341 48557 7362 48613
rect 7264 48536 7362 48557
rect 7660 48613 7758 48634
rect 7660 48557 7681 48613
rect 7737 48557 7758 48613
rect 7660 48536 7758 48557
rect 6025 48262 6123 48283
rect 6025 48206 6046 48262
rect 6102 48206 6123 48262
rect 6025 48185 6123 48206
rect 6450 48204 6548 48225
rect 6450 48148 6471 48204
rect 6527 48148 6548 48204
rect 6450 48127 6548 48148
rect 6882 48204 6980 48225
rect 6882 48148 6903 48204
rect 6959 48148 6980 48204
rect 6882 48127 6980 48148
rect 7264 48218 7362 48239
rect 7264 48162 7285 48218
rect 7341 48162 7362 48218
rect 7264 48141 7362 48162
rect 7660 48218 7758 48239
rect 7660 48162 7681 48218
rect 7737 48162 7758 48218
rect 7660 48141 7758 48162
rect 6025 47846 6123 47867
rect 6025 47790 6046 47846
rect 6102 47790 6123 47846
rect 6025 47769 6123 47790
rect 6450 47846 6548 47867
rect 6450 47790 6471 47846
rect 6527 47790 6548 47846
rect 6450 47769 6548 47790
rect 6882 47846 6980 47867
rect 6882 47790 6903 47846
rect 6959 47790 6980 47846
rect 6882 47769 6980 47790
rect 7264 47823 7362 47844
rect 7264 47767 7285 47823
rect 7341 47767 7362 47823
rect 7264 47746 7362 47767
rect 7660 47823 7758 47844
rect 7660 47767 7681 47823
rect 7737 47767 7758 47823
rect 7660 47746 7758 47767
rect 6025 47472 6123 47493
rect 6025 47416 6046 47472
rect 6102 47416 6123 47472
rect 6025 47395 6123 47416
rect 6450 47414 6548 47435
rect 6450 47358 6471 47414
rect 6527 47358 6548 47414
rect 6450 47337 6548 47358
rect 6882 47414 6980 47435
rect 6882 47358 6903 47414
rect 6959 47358 6980 47414
rect 6882 47337 6980 47358
rect 7264 47428 7362 47449
rect 7264 47372 7285 47428
rect 7341 47372 7362 47428
rect 7264 47351 7362 47372
rect 7660 47428 7758 47449
rect 7660 47372 7681 47428
rect 7737 47372 7758 47428
rect 7660 47351 7758 47372
rect 6025 47056 6123 47077
rect 6025 47000 6046 47056
rect 6102 47000 6123 47056
rect 6025 46979 6123 47000
rect 6450 47056 6548 47077
rect 6450 47000 6471 47056
rect 6527 47000 6548 47056
rect 6450 46979 6548 47000
rect 6882 47056 6980 47077
rect 6882 47000 6903 47056
rect 6959 47000 6980 47056
rect 6882 46979 6980 47000
rect 7264 47033 7362 47054
rect 7264 46977 7285 47033
rect 7341 46977 7362 47033
rect 7264 46956 7362 46977
rect 7660 47033 7758 47054
rect 7660 46977 7681 47033
rect 7737 46977 7758 47033
rect 7660 46956 7758 46977
rect 6025 46682 6123 46703
rect 6025 46626 6046 46682
rect 6102 46626 6123 46682
rect 6025 46605 6123 46626
rect 6450 46624 6548 46645
rect 6450 46568 6471 46624
rect 6527 46568 6548 46624
rect 6450 46547 6548 46568
rect 6882 46624 6980 46645
rect 6882 46568 6903 46624
rect 6959 46568 6980 46624
rect 6882 46547 6980 46568
rect 7264 46638 7362 46659
rect 7264 46582 7285 46638
rect 7341 46582 7362 46638
rect 7264 46561 7362 46582
rect 7660 46638 7758 46659
rect 7660 46582 7681 46638
rect 7737 46582 7758 46638
rect 7660 46561 7758 46582
rect 6025 46266 6123 46287
rect 6025 46210 6046 46266
rect 6102 46210 6123 46266
rect 6025 46189 6123 46210
rect 6450 46266 6548 46287
rect 6450 46210 6471 46266
rect 6527 46210 6548 46266
rect 6450 46189 6548 46210
rect 6882 46266 6980 46287
rect 6882 46210 6903 46266
rect 6959 46210 6980 46266
rect 6882 46189 6980 46210
rect 7264 46243 7362 46264
rect 7264 46187 7285 46243
rect 7341 46187 7362 46243
rect 7264 46166 7362 46187
rect 7660 46243 7758 46264
rect 7660 46187 7681 46243
rect 7737 46187 7758 46243
rect 7660 46166 7758 46187
rect 6025 45892 6123 45913
rect 6025 45836 6046 45892
rect 6102 45836 6123 45892
rect 6025 45815 6123 45836
rect 6450 45834 6548 45855
rect 6450 45778 6471 45834
rect 6527 45778 6548 45834
rect 6450 45757 6548 45778
rect 6882 45834 6980 45855
rect 6882 45778 6903 45834
rect 6959 45778 6980 45834
rect 6882 45757 6980 45778
rect 7264 45848 7362 45869
rect 7264 45792 7285 45848
rect 7341 45792 7362 45848
rect 7264 45771 7362 45792
rect 7660 45848 7758 45869
rect 7660 45792 7681 45848
rect 7737 45792 7758 45848
rect 7660 45771 7758 45792
rect 6025 45476 6123 45497
rect 6025 45420 6046 45476
rect 6102 45420 6123 45476
rect 6025 45399 6123 45420
rect 6450 45476 6548 45497
rect 6450 45420 6471 45476
rect 6527 45420 6548 45476
rect 6450 45399 6548 45420
rect 6882 45476 6980 45497
rect 6882 45420 6903 45476
rect 6959 45420 6980 45476
rect 6882 45399 6980 45420
rect 7264 45453 7362 45474
rect 7264 45397 7285 45453
rect 7341 45397 7362 45453
rect 7264 45376 7362 45397
rect 7660 45453 7758 45474
rect 7660 45397 7681 45453
rect 7737 45397 7758 45453
rect 7660 45376 7758 45397
rect 6025 45102 6123 45123
rect 6025 45046 6046 45102
rect 6102 45046 6123 45102
rect 6025 45025 6123 45046
rect 6450 45044 6548 45065
rect 6450 44988 6471 45044
rect 6527 44988 6548 45044
rect 6450 44967 6548 44988
rect 6882 45044 6980 45065
rect 6882 44988 6903 45044
rect 6959 44988 6980 45044
rect 6882 44967 6980 44988
rect 7264 45058 7362 45079
rect 7264 45002 7285 45058
rect 7341 45002 7362 45058
rect 7264 44981 7362 45002
rect 7660 45058 7758 45079
rect 7660 45002 7681 45058
rect 7737 45002 7758 45058
rect 7660 44981 7758 45002
rect 6025 44686 6123 44707
rect 6025 44630 6046 44686
rect 6102 44630 6123 44686
rect 6025 44609 6123 44630
rect 6450 44686 6548 44707
rect 6450 44630 6471 44686
rect 6527 44630 6548 44686
rect 6450 44609 6548 44630
rect 6882 44686 6980 44707
rect 6882 44630 6903 44686
rect 6959 44630 6980 44686
rect 6882 44609 6980 44630
rect 7264 44663 7362 44684
rect 7264 44607 7285 44663
rect 7341 44607 7362 44663
rect 7264 44586 7362 44607
rect 7660 44663 7758 44684
rect 7660 44607 7681 44663
rect 7737 44607 7758 44663
rect 7660 44586 7758 44607
rect 6025 44312 6123 44333
rect 6025 44256 6046 44312
rect 6102 44256 6123 44312
rect 6025 44235 6123 44256
rect 6450 44254 6548 44275
rect 6450 44198 6471 44254
rect 6527 44198 6548 44254
rect 6450 44177 6548 44198
rect 6882 44254 6980 44275
rect 6882 44198 6903 44254
rect 6959 44198 6980 44254
rect 6882 44177 6980 44198
rect 7264 44268 7362 44289
rect 7264 44212 7285 44268
rect 7341 44212 7362 44268
rect 7264 44191 7362 44212
rect 7660 44268 7758 44289
rect 7660 44212 7681 44268
rect 7737 44212 7758 44268
rect 7660 44191 7758 44212
rect 6025 43896 6123 43917
rect 6025 43840 6046 43896
rect 6102 43840 6123 43896
rect 6025 43819 6123 43840
rect 6450 43896 6548 43917
rect 6450 43840 6471 43896
rect 6527 43840 6548 43896
rect 6450 43819 6548 43840
rect 6882 43896 6980 43917
rect 6882 43840 6903 43896
rect 6959 43840 6980 43896
rect 6882 43819 6980 43840
rect 7264 43873 7362 43894
rect 7264 43817 7285 43873
rect 7341 43817 7362 43873
rect 7264 43796 7362 43817
rect 7660 43873 7758 43894
rect 7660 43817 7681 43873
rect 7737 43817 7758 43873
rect 7660 43796 7758 43817
rect 6025 43522 6123 43543
rect 6025 43466 6046 43522
rect 6102 43466 6123 43522
rect 6025 43445 6123 43466
rect 6450 43464 6548 43485
rect 6450 43408 6471 43464
rect 6527 43408 6548 43464
rect 6450 43387 6548 43408
rect 6882 43464 6980 43485
rect 6882 43408 6903 43464
rect 6959 43408 6980 43464
rect 6882 43387 6980 43408
rect 7264 43478 7362 43499
rect 7264 43422 7285 43478
rect 7341 43422 7362 43478
rect 7264 43401 7362 43422
rect 7660 43478 7758 43499
rect 7660 43422 7681 43478
rect 7737 43422 7758 43478
rect 7660 43401 7758 43422
rect 6025 43106 6123 43127
rect 6025 43050 6046 43106
rect 6102 43050 6123 43106
rect 6025 43029 6123 43050
rect 6450 43106 6548 43127
rect 6450 43050 6471 43106
rect 6527 43050 6548 43106
rect 6450 43029 6548 43050
rect 6882 43106 6980 43127
rect 6882 43050 6903 43106
rect 6959 43050 6980 43106
rect 6882 43029 6980 43050
rect 7264 43083 7362 43104
rect 7264 43027 7285 43083
rect 7341 43027 7362 43083
rect 7264 43006 7362 43027
rect 7660 43083 7758 43104
rect 7660 43027 7681 43083
rect 7737 43027 7758 43083
rect 7660 43006 7758 43027
rect 6025 42732 6123 42753
rect 6025 42676 6046 42732
rect 6102 42676 6123 42732
rect 6025 42655 6123 42676
rect 6450 42674 6548 42695
rect 6450 42618 6471 42674
rect 6527 42618 6548 42674
rect 6450 42597 6548 42618
rect 6882 42674 6980 42695
rect 6882 42618 6903 42674
rect 6959 42618 6980 42674
rect 6882 42597 6980 42618
rect 7264 42688 7362 42709
rect 7264 42632 7285 42688
rect 7341 42632 7362 42688
rect 7264 42611 7362 42632
rect 7660 42688 7758 42709
rect 7660 42632 7681 42688
rect 7737 42632 7758 42688
rect 7660 42611 7758 42632
rect 6025 42316 6123 42337
rect 6025 42260 6046 42316
rect 6102 42260 6123 42316
rect 6025 42239 6123 42260
rect 6450 42316 6548 42337
rect 6450 42260 6471 42316
rect 6527 42260 6548 42316
rect 6450 42239 6548 42260
rect 6882 42316 6980 42337
rect 6882 42260 6903 42316
rect 6959 42260 6980 42316
rect 6882 42239 6980 42260
rect 7264 42293 7362 42314
rect 7264 42237 7285 42293
rect 7341 42237 7362 42293
rect 7264 42216 7362 42237
rect 7660 42293 7758 42314
rect 7660 42237 7681 42293
rect 7737 42237 7758 42293
rect 7660 42216 7758 42237
rect 6025 41942 6123 41963
rect 6025 41886 6046 41942
rect 6102 41886 6123 41942
rect 6025 41865 6123 41886
rect 6450 41884 6548 41905
rect 6450 41828 6471 41884
rect 6527 41828 6548 41884
rect 6450 41807 6548 41828
rect 6882 41884 6980 41905
rect 6882 41828 6903 41884
rect 6959 41828 6980 41884
rect 6882 41807 6980 41828
rect 7264 41898 7362 41919
rect 7264 41842 7285 41898
rect 7341 41842 7362 41898
rect 7264 41821 7362 41842
rect 7660 41898 7758 41919
rect 7660 41842 7681 41898
rect 7737 41842 7758 41898
rect 7660 41821 7758 41842
rect 6025 41526 6123 41547
rect 6025 41470 6046 41526
rect 6102 41470 6123 41526
rect 6025 41449 6123 41470
rect 6450 41526 6548 41547
rect 6450 41470 6471 41526
rect 6527 41470 6548 41526
rect 6450 41449 6548 41470
rect 6882 41526 6980 41547
rect 6882 41470 6903 41526
rect 6959 41470 6980 41526
rect 6882 41449 6980 41470
rect 7264 41503 7362 41524
rect 7264 41447 7285 41503
rect 7341 41447 7362 41503
rect 7264 41426 7362 41447
rect 7660 41503 7758 41524
rect 7660 41447 7681 41503
rect 7737 41447 7758 41503
rect 7660 41426 7758 41447
rect 6025 41152 6123 41173
rect 6025 41096 6046 41152
rect 6102 41096 6123 41152
rect 6025 41075 6123 41096
rect 6450 41094 6548 41115
rect 6450 41038 6471 41094
rect 6527 41038 6548 41094
rect 6450 41017 6548 41038
rect 6882 41094 6980 41115
rect 6882 41038 6903 41094
rect 6959 41038 6980 41094
rect 6882 41017 6980 41038
rect 7264 41108 7362 41129
rect 7264 41052 7285 41108
rect 7341 41052 7362 41108
rect 7264 41031 7362 41052
rect 7660 41108 7758 41129
rect 7660 41052 7681 41108
rect 7737 41052 7758 41108
rect 7660 41031 7758 41052
rect 6025 40736 6123 40757
rect 6025 40680 6046 40736
rect 6102 40680 6123 40736
rect 6025 40659 6123 40680
rect 6450 40736 6548 40757
rect 6450 40680 6471 40736
rect 6527 40680 6548 40736
rect 6450 40659 6548 40680
rect 6882 40736 6980 40757
rect 6882 40680 6903 40736
rect 6959 40680 6980 40736
rect 6882 40659 6980 40680
rect 7264 40713 7362 40734
rect 7264 40657 7285 40713
rect 7341 40657 7362 40713
rect 7264 40636 7362 40657
rect 7660 40713 7758 40734
rect 7660 40657 7681 40713
rect 7737 40657 7758 40713
rect 7660 40636 7758 40657
rect 6025 40362 6123 40383
rect 6025 40306 6046 40362
rect 6102 40306 6123 40362
rect 6025 40285 6123 40306
rect 6450 40304 6548 40325
rect 6450 40248 6471 40304
rect 6527 40248 6548 40304
rect 6450 40227 6548 40248
rect 6882 40304 6980 40325
rect 6882 40248 6903 40304
rect 6959 40248 6980 40304
rect 6882 40227 6980 40248
rect 7264 40318 7362 40339
rect 7264 40262 7285 40318
rect 7341 40262 7362 40318
rect 7264 40241 7362 40262
rect 7660 40318 7758 40339
rect 7660 40262 7681 40318
rect 7737 40262 7758 40318
rect 7660 40241 7758 40262
rect 6025 39946 6123 39967
rect 6025 39890 6046 39946
rect 6102 39890 6123 39946
rect 6025 39869 6123 39890
rect 6450 39946 6548 39967
rect 6450 39890 6471 39946
rect 6527 39890 6548 39946
rect 6450 39869 6548 39890
rect 6882 39946 6980 39967
rect 6882 39890 6903 39946
rect 6959 39890 6980 39946
rect 6882 39869 6980 39890
rect 7264 39923 7362 39944
rect 7264 39867 7285 39923
rect 7341 39867 7362 39923
rect 7264 39846 7362 39867
rect 7660 39923 7758 39944
rect 7660 39867 7681 39923
rect 7737 39867 7758 39923
rect 7660 39846 7758 39867
rect 6025 39572 6123 39593
rect 6025 39516 6046 39572
rect 6102 39516 6123 39572
rect 6025 39495 6123 39516
rect 6450 39514 6548 39535
rect 6450 39458 6471 39514
rect 6527 39458 6548 39514
rect 6450 39437 6548 39458
rect 6882 39514 6980 39535
rect 6882 39458 6903 39514
rect 6959 39458 6980 39514
rect 6882 39437 6980 39458
rect 7264 39528 7362 39549
rect 7264 39472 7285 39528
rect 7341 39472 7362 39528
rect 7264 39451 7362 39472
rect 7660 39528 7758 39549
rect 7660 39472 7681 39528
rect 7737 39472 7758 39528
rect 7660 39451 7758 39472
rect 6025 39156 6123 39177
rect 6025 39100 6046 39156
rect 6102 39100 6123 39156
rect 6025 39079 6123 39100
rect 6450 39156 6548 39177
rect 6450 39100 6471 39156
rect 6527 39100 6548 39156
rect 6450 39079 6548 39100
rect 6882 39156 6980 39177
rect 6882 39100 6903 39156
rect 6959 39100 6980 39156
rect 6882 39079 6980 39100
rect 7264 39133 7362 39154
rect 7264 39077 7285 39133
rect 7341 39077 7362 39133
rect 7264 39056 7362 39077
rect 7660 39133 7758 39154
rect 7660 39077 7681 39133
rect 7737 39077 7758 39133
rect 7660 39056 7758 39077
rect 6025 38782 6123 38803
rect 6025 38726 6046 38782
rect 6102 38726 6123 38782
rect 6025 38705 6123 38726
rect 6450 38724 6548 38745
rect 6450 38668 6471 38724
rect 6527 38668 6548 38724
rect 6450 38647 6548 38668
rect 6882 38724 6980 38745
rect 6882 38668 6903 38724
rect 6959 38668 6980 38724
rect 6882 38647 6980 38668
rect 7264 38738 7362 38759
rect 7264 38682 7285 38738
rect 7341 38682 7362 38738
rect 7264 38661 7362 38682
rect 7660 38738 7758 38759
rect 7660 38682 7681 38738
rect 7737 38682 7758 38738
rect 7660 38661 7758 38682
rect 6025 38366 6123 38387
rect 6025 38310 6046 38366
rect 6102 38310 6123 38366
rect 6025 38289 6123 38310
rect 6450 38366 6548 38387
rect 6450 38310 6471 38366
rect 6527 38310 6548 38366
rect 6450 38289 6548 38310
rect 6882 38366 6980 38387
rect 6882 38310 6903 38366
rect 6959 38310 6980 38366
rect 6882 38289 6980 38310
rect 7264 38343 7362 38364
rect 7264 38287 7285 38343
rect 7341 38287 7362 38343
rect 7264 38266 7362 38287
rect 7660 38343 7758 38364
rect 7660 38287 7681 38343
rect 7737 38287 7758 38343
rect 7660 38266 7758 38287
rect 6025 37992 6123 38013
rect 6025 37936 6046 37992
rect 6102 37936 6123 37992
rect 6025 37915 6123 37936
rect 6450 37934 6548 37955
rect 6450 37878 6471 37934
rect 6527 37878 6548 37934
rect 6450 37857 6548 37878
rect 6882 37934 6980 37955
rect 6882 37878 6903 37934
rect 6959 37878 6980 37934
rect 6882 37857 6980 37878
rect 7264 37948 7362 37969
rect 7264 37892 7285 37948
rect 7341 37892 7362 37948
rect 7264 37871 7362 37892
rect 7660 37948 7758 37969
rect 7660 37892 7681 37948
rect 7737 37892 7758 37948
rect 7660 37871 7758 37892
rect 6025 37576 6123 37597
rect 6025 37520 6046 37576
rect 6102 37520 6123 37576
rect 6025 37499 6123 37520
rect 6450 37576 6548 37597
rect 6450 37520 6471 37576
rect 6527 37520 6548 37576
rect 6450 37499 6548 37520
rect 6882 37576 6980 37597
rect 6882 37520 6903 37576
rect 6959 37520 6980 37576
rect 6882 37499 6980 37520
rect 7264 37553 7362 37574
rect 7264 37497 7285 37553
rect 7341 37497 7362 37553
rect 7264 37476 7362 37497
rect 7660 37553 7758 37574
rect 7660 37497 7681 37553
rect 7737 37497 7758 37553
rect 7660 37476 7758 37497
rect 6025 37202 6123 37223
rect 6025 37146 6046 37202
rect 6102 37146 6123 37202
rect 6025 37125 6123 37146
rect 6450 37144 6548 37165
rect 6450 37088 6471 37144
rect 6527 37088 6548 37144
rect 6450 37067 6548 37088
rect 6882 37144 6980 37165
rect 6882 37088 6903 37144
rect 6959 37088 6980 37144
rect 6882 37067 6980 37088
rect 7264 37158 7362 37179
rect 7264 37102 7285 37158
rect 7341 37102 7362 37158
rect 7264 37081 7362 37102
rect 7660 37158 7758 37179
rect 7660 37102 7681 37158
rect 7737 37102 7758 37158
rect 7660 37081 7758 37102
rect 6025 36786 6123 36807
rect 6025 36730 6046 36786
rect 6102 36730 6123 36786
rect 6025 36709 6123 36730
rect 6450 36786 6548 36807
rect 6450 36730 6471 36786
rect 6527 36730 6548 36786
rect 6450 36709 6548 36730
rect 6882 36786 6980 36807
rect 6882 36730 6903 36786
rect 6959 36730 6980 36786
rect 6882 36709 6980 36730
rect 7264 36763 7362 36784
rect 7264 36707 7285 36763
rect 7341 36707 7362 36763
rect 7264 36686 7362 36707
rect 7660 36763 7758 36784
rect 7660 36707 7681 36763
rect 7737 36707 7758 36763
rect 7660 36686 7758 36707
rect 6025 36412 6123 36433
rect 6025 36356 6046 36412
rect 6102 36356 6123 36412
rect 6025 36335 6123 36356
rect 6450 36354 6548 36375
rect 6450 36298 6471 36354
rect 6527 36298 6548 36354
rect 6450 36277 6548 36298
rect 6882 36354 6980 36375
rect 6882 36298 6903 36354
rect 6959 36298 6980 36354
rect 6882 36277 6980 36298
rect 7264 36368 7362 36389
rect 7264 36312 7285 36368
rect 7341 36312 7362 36368
rect 7264 36291 7362 36312
rect 7660 36368 7758 36389
rect 7660 36312 7681 36368
rect 7737 36312 7758 36368
rect 7660 36291 7758 36312
rect 6025 35996 6123 36017
rect 6025 35940 6046 35996
rect 6102 35940 6123 35996
rect 6025 35919 6123 35940
rect 6450 35996 6548 36017
rect 6450 35940 6471 35996
rect 6527 35940 6548 35996
rect 6450 35919 6548 35940
rect 6882 35996 6980 36017
rect 6882 35940 6903 35996
rect 6959 35940 6980 35996
rect 6882 35919 6980 35940
rect 7264 35973 7362 35994
rect 7264 35917 7285 35973
rect 7341 35917 7362 35973
rect 7264 35896 7362 35917
rect 7660 35973 7758 35994
rect 7660 35917 7681 35973
rect 7737 35917 7758 35973
rect 7660 35896 7758 35917
rect 6025 35622 6123 35643
rect 6025 35566 6046 35622
rect 6102 35566 6123 35622
rect 6025 35545 6123 35566
rect 6450 35564 6548 35585
rect 6450 35508 6471 35564
rect 6527 35508 6548 35564
rect 6450 35487 6548 35508
rect 6882 35564 6980 35585
rect 6882 35508 6903 35564
rect 6959 35508 6980 35564
rect 6882 35487 6980 35508
rect 7264 35578 7362 35599
rect 7264 35522 7285 35578
rect 7341 35522 7362 35578
rect 7264 35501 7362 35522
rect 7660 35578 7758 35599
rect 7660 35522 7681 35578
rect 7737 35522 7758 35578
rect 7660 35501 7758 35522
rect 6025 35206 6123 35227
rect 6025 35150 6046 35206
rect 6102 35150 6123 35206
rect 6025 35129 6123 35150
rect 6450 35206 6548 35227
rect 6450 35150 6471 35206
rect 6527 35150 6548 35206
rect 6450 35129 6548 35150
rect 6882 35206 6980 35227
rect 6882 35150 6903 35206
rect 6959 35150 6980 35206
rect 6882 35129 6980 35150
rect 7264 35183 7362 35204
rect 7264 35127 7285 35183
rect 7341 35127 7362 35183
rect 7264 35106 7362 35127
rect 7660 35183 7758 35204
rect 7660 35127 7681 35183
rect 7737 35127 7758 35183
rect 7660 35106 7758 35127
rect 6025 34832 6123 34853
rect 6025 34776 6046 34832
rect 6102 34776 6123 34832
rect 6025 34755 6123 34776
rect 6450 34774 6548 34795
rect 6450 34718 6471 34774
rect 6527 34718 6548 34774
rect 6450 34697 6548 34718
rect 6882 34774 6980 34795
rect 6882 34718 6903 34774
rect 6959 34718 6980 34774
rect 6882 34697 6980 34718
rect 7264 34788 7362 34809
rect 7264 34732 7285 34788
rect 7341 34732 7362 34788
rect 7264 34711 7362 34732
rect 7660 34788 7758 34809
rect 7660 34732 7681 34788
rect 7737 34732 7758 34788
rect 7660 34711 7758 34732
rect 6025 34416 6123 34437
rect 6025 34360 6046 34416
rect 6102 34360 6123 34416
rect 6025 34339 6123 34360
rect 6450 34416 6548 34437
rect 6450 34360 6471 34416
rect 6527 34360 6548 34416
rect 6450 34339 6548 34360
rect 6882 34416 6980 34437
rect 6882 34360 6903 34416
rect 6959 34360 6980 34416
rect 6882 34339 6980 34360
rect 7264 34393 7362 34414
rect 7264 34337 7285 34393
rect 7341 34337 7362 34393
rect 7264 34316 7362 34337
rect 7660 34393 7758 34414
rect 7660 34337 7681 34393
rect 7737 34337 7758 34393
rect 7660 34316 7758 34337
rect 6025 34042 6123 34063
rect 6025 33986 6046 34042
rect 6102 33986 6123 34042
rect 6025 33965 6123 33986
rect 6450 33984 6548 34005
rect 6450 33928 6471 33984
rect 6527 33928 6548 33984
rect 6450 33907 6548 33928
rect 6882 33984 6980 34005
rect 6882 33928 6903 33984
rect 6959 33928 6980 33984
rect 6882 33907 6980 33928
rect 7264 33998 7362 34019
rect 7264 33942 7285 33998
rect 7341 33942 7362 33998
rect 7264 33921 7362 33942
rect 7660 33998 7758 34019
rect 7660 33942 7681 33998
rect 7737 33942 7758 33998
rect 7660 33921 7758 33942
rect 6025 33626 6123 33647
rect 6025 33570 6046 33626
rect 6102 33570 6123 33626
rect 6025 33549 6123 33570
rect 6450 33626 6548 33647
rect 6450 33570 6471 33626
rect 6527 33570 6548 33626
rect 6450 33549 6548 33570
rect 6882 33626 6980 33647
rect 6882 33570 6903 33626
rect 6959 33570 6980 33626
rect 6882 33549 6980 33570
rect 7264 33603 7362 33624
rect 7264 33547 7285 33603
rect 7341 33547 7362 33603
rect 7264 33526 7362 33547
rect 7660 33603 7758 33624
rect 7660 33547 7681 33603
rect 7737 33547 7758 33603
rect 7660 33526 7758 33547
rect 6025 33252 6123 33273
rect 6025 33196 6046 33252
rect 6102 33196 6123 33252
rect 6025 33175 6123 33196
rect 6450 33194 6548 33215
rect 6450 33138 6471 33194
rect 6527 33138 6548 33194
rect 6450 33117 6548 33138
rect 6882 33194 6980 33215
rect 6882 33138 6903 33194
rect 6959 33138 6980 33194
rect 6882 33117 6980 33138
rect 7264 33208 7362 33229
rect 7264 33152 7285 33208
rect 7341 33152 7362 33208
rect 7264 33131 7362 33152
rect 7660 33208 7758 33229
rect 7660 33152 7681 33208
rect 7737 33152 7758 33208
rect 7660 33131 7758 33152
rect 6025 32836 6123 32857
rect 6025 32780 6046 32836
rect 6102 32780 6123 32836
rect 6025 32759 6123 32780
rect 6450 32836 6548 32857
rect 6450 32780 6471 32836
rect 6527 32780 6548 32836
rect 6450 32759 6548 32780
rect 6882 32836 6980 32857
rect 6882 32780 6903 32836
rect 6959 32780 6980 32836
rect 6882 32759 6980 32780
rect 7264 32813 7362 32834
rect 7264 32757 7285 32813
rect 7341 32757 7362 32813
rect 7264 32736 7362 32757
rect 7660 32813 7758 32834
rect 7660 32757 7681 32813
rect 7737 32757 7758 32813
rect 7660 32736 7758 32757
rect 6025 32462 6123 32483
rect 6025 32406 6046 32462
rect 6102 32406 6123 32462
rect 6025 32385 6123 32406
rect 6450 32404 6548 32425
rect 6450 32348 6471 32404
rect 6527 32348 6548 32404
rect 6450 32327 6548 32348
rect 6882 32404 6980 32425
rect 6882 32348 6903 32404
rect 6959 32348 6980 32404
rect 6882 32327 6980 32348
rect 7264 32418 7362 32439
rect 7264 32362 7285 32418
rect 7341 32362 7362 32418
rect 7264 32341 7362 32362
rect 7660 32418 7758 32439
rect 7660 32362 7681 32418
rect 7737 32362 7758 32418
rect 7660 32341 7758 32362
rect 6025 32046 6123 32067
rect 6025 31990 6046 32046
rect 6102 31990 6123 32046
rect 6025 31969 6123 31990
rect 6450 32046 6548 32067
rect 6450 31990 6471 32046
rect 6527 31990 6548 32046
rect 6450 31969 6548 31990
rect 6882 32046 6980 32067
rect 6882 31990 6903 32046
rect 6959 31990 6980 32046
rect 6882 31969 6980 31990
rect 7264 32023 7362 32044
rect 7264 31967 7285 32023
rect 7341 31967 7362 32023
rect 7264 31946 7362 31967
rect 7660 32023 7758 32044
rect 7660 31967 7681 32023
rect 7737 31967 7758 32023
rect 7660 31946 7758 31967
rect 6025 31672 6123 31693
rect 6025 31616 6046 31672
rect 6102 31616 6123 31672
rect 6025 31595 6123 31616
rect 6450 31614 6548 31635
rect 6450 31558 6471 31614
rect 6527 31558 6548 31614
rect 6450 31537 6548 31558
rect 6882 31614 6980 31635
rect 6882 31558 6903 31614
rect 6959 31558 6980 31614
rect 6882 31537 6980 31558
rect 7264 31628 7362 31649
rect 7264 31572 7285 31628
rect 7341 31572 7362 31628
rect 7264 31551 7362 31572
rect 7660 31628 7758 31649
rect 7660 31572 7681 31628
rect 7737 31572 7758 31628
rect 7660 31551 7758 31572
rect 6025 31256 6123 31277
rect 6025 31200 6046 31256
rect 6102 31200 6123 31256
rect 6025 31179 6123 31200
rect 6450 31256 6548 31277
rect 6450 31200 6471 31256
rect 6527 31200 6548 31256
rect 6450 31179 6548 31200
rect 6882 31256 6980 31277
rect 6882 31200 6903 31256
rect 6959 31200 6980 31256
rect 6882 31179 6980 31200
rect 7264 31233 7362 31254
rect 7264 31177 7285 31233
rect 7341 31177 7362 31233
rect 7264 31156 7362 31177
rect 7660 31233 7758 31254
rect 7660 31177 7681 31233
rect 7737 31177 7758 31233
rect 7660 31156 7758 31177
rect 6025 30882 6123 30903
rect 6025 30826 6046 30882
rect 6102 30826 6123 30882
rect 6025 30805 6123 30826
rect 6450 30824 6548 30845
rect 6450 30768 6471 30824
rect 6527 30768 6548 30824
rect 6450 30747 6548 30768
rect 6882 30824 6980 30845
rect 6882 30768 6903 30824
rect 6959 30768 6980 30824
rect 6882 30747 6980 30768
rect 7264 30838 7362 30859
rect 7264 30782 7285 30838
rect 7341 30782 7362 30838
rect 7264 30761 7362 30782
rect 7660 30838 7758 30859
rect 7660 30782 7681 30838
rect 7737 30782 7758 30838
rect 7660 30761 7758 30782
rect 6025 30466 6123 30487
rect 6025 30410 6046 30466
rect 6102 30410 6123 30466
rect 6025 30389 6123 30410
rect 6450 30466 6548 30487
rect 6450 30410 6471 30466
rect 6527 30410 6548 30466
rect 6450 30389 6548 30410
rect 6882 30466 6980 30487
rect 6882 30410 6903 30466
rect 6959 30410 6980 30466
rect 6882 30389 6980 30410
rect 7264 30443 7362 30464
rect 7264 30387 7285 30443
rect 7341 30387 7362 30443
rect 7264 30366 7362 30387
rect 7660 30443 7758 30464
rect 7660 30387 7681 30443
rect 7737 30387 7758 30443
rect 7660 30366 7758 30387
rect 6025 30092 6123 30113
rect 6025 30036 6046 30092
rect 6102 30036 6123 30092
rect 6025 30015 6123 30036
rect 6450 30034 6548 30055
rect 6450 29978 6471 30034
rect 6527 29978 6548 30034
rect 6450 29957 6548 29978
rect 6882 30034 6980 30055
rect 6882 29978 6903 30034
rect 6959 29978 6980 30034
rect 6882 29957 6980 29978
rect 7264 30048 7362 30069
rect 7264 29992 7285 30048
rect 7341 29992 7362 30048
rect 7264 29971 7362 29992
rect 7660 30048 7758 30069
rect 7660 29992 7681 30048
rect 7737 29992 7758 30048
rect 7660 29971 7758 29992
rect 6025 29676 6123 29697
rect 6025 29620 6046 29676
rect 6102 29620 6123 29676
rect 6025 29599 6123 29620
rect 6450 29676 6548 29697
rect 6450 29620 6471 29676
rect 6527 29620 6548 29676
rect 6450 29599 6548 29620
rect 6882 29676 6980 29697
rect 6882 29620 6903 29676
rect 6959 29620 6980 29676
rect 6882 29599 6980 29620
rect 7264 29653 7362 29674
rect 7264 29597 7285 29653
rect 7341 29597 7362 29653
rect 7264 29576 7362 29597
rect 7660 29653 7758 29674
rect 7660 29597 7681 29653
rect 7737 29597 7758 29653
rect 7660 29576 7758 29597
rect 6025 29302 6123 29323
rect 6025 29246 6046 29302
rect 6102 29246 6123 29302
rect 6025 29225 6123 29246
rect 6450 29244 6548 29265
rect 6450 29188 6471 29244
rect 6527 29188 6548 29244
rect 6450 29167 6548 29188
rect 6882 29244 6980 29265
rect 6882 29188 6903 29244
rect 6959 29188 6980 29244
rect 6882 29167 6980 29188
rect 7264 29258 7362 29279
rect 7264 29202 7285 29258
rect 7341 29202 7362 29258
rect 7264 29181 7362 29202
rect 7660 29258 7758 29279
rect 7660 29202 7681 29258
rect 7737 29202 7758 29258
rect 7660 29181 7758 29202
rect 6025 28886 6123 28907
rect 6025 28830 6046 28886
rect 6102 28830 6123 28886
rect 6025 28809 6123 28830
rect 6450 28886 6548 28907
rect 6450 28830 6471 28886
rect 6527 28830 6548 28886
rect 6450 28809 6548 28830
rect 6882 28886 6980 28907
rect 6882 28830 6903 28886
rect 6959 28830 6980 28886
rect 6882 28809 6980 28830
rect 7264 28863 7362 28884
rect 7264 28807 7285 28863
rect 7341 28807 7362 28863
rect 7264 28786 7362 28807
rect 7660 28863 7758 28884
rect 7660 28807 7681 28863
rect 7737 28807 7758 28863
rect 7660 28786 7758 28807
rect 6025 28512 6123 28533
rect 6025 28456 6046 28512
rect 6102 28456 6123 28512
rect 6025 28435 6123 28456
rect 6450 28454 6548 28475
rect 6450 28398 6471 28454
rect 6527 28398 6548 28454
rect 6450 28377 6548 28398
rect 6882 28454 6980 28475
rect 6882 28398 6903 28454
rect 6959 28398 6980 28454
rect 6882 28377 6980 28398
rect 7264 28468 7362 28489
rect 7264 28412 7285 28468
rect 7341 28412 7362 28468
rect 7264 28391 7362 28412
rect 7660 28468 7758 28489
rect 7660 28412 7681 28468
rect 7737 28412 7758 28468
rect 7660 28391 7758 28412
rect 6025 28096 6123 28117
rect 6025 28040 6046 28096
rect 6102 28040 6123 28096
rect 6025 28019 6123 28040
rect 6450 28096 6548 28117
rect 6450 28040 6471 28096
rect 6527 28040 6548 28096
rect 6450 28019 6548 28040
rect 6882 28096 6980 28117
rect 6882 28040 6903 28096
rect 6959 28040 6980 28096
rect 6882 28019 6980 28040
rect 7264 28073 7362 28094
rect 7264 28017 7285 28073
rect 7341 28017 7362 28073
rect 7264 27996 7362 28017
rect 7660 28073 7758 28094
rect 7660 28017 7681 28073
rect 7737 28017 7758 28073
rect 7660 27996 7758 28017
rect 6025 27722 6123 27743
rect 6025 27666 6046 27722
rect 6102 27666 6123 27722
rect 6025 27645 6123 27666
rect 6450 27664 6548 27685
rect 6450 27608 6471 27664
rect 6527 27608 6548 27664
rect 6450 27587 6548 27608
rect 6882 27664 6980 27685
rect 6882 27608 6903 27664
rect 6959 27608 6980 27664
rect 6882 27587 6980 27608
rect 7264 27678 7362 27699
rect 7264 27622 7285 27678
rect 7341 27622 7362 27678
rect 7264 27601 7362 27622
rect 7660 27678 7758 27699
rect 7660 27622 7681 27678
rect 7737 27622 7758 27678
rect 7660 27601 7758 27622
rect 6025 27306 6123 27327
rect 6025 27250 6046 27306
rect 6102 27250 6123 27306
rect 6025 27229 6123 27250
rect 6450 27306 6548 27327
rect 6450 27250 6471 27306
rect 6527 27250 6548 27306
rect 6450 27229 6548 27250
rect 6882 27306 6980 27327
rect 6882 27250 6903 27306
rect 6959 27250 6980 27306
rect 6882 27229 6980 27250
rect 7264 27283 7362 27304
rect 7264 27227 7285 27283
rect 7341 27227 7362 27283
rect 7264 27206 7362 27227
rect 7660 27283 7758 27304
rect 7660 27227 7681 27283
rect 7737 27227 7758 27283
rect 7660 27206 7758 27227
rect 6025 26932 6123 26953
rect 6025 26876 6046 26932
rect 6102 26876 6123 26932
rect 6025 26855 6123 26876
rect 6450 26874 6548 26895
rect 6450 26818 6471 26874
rect 6527 26818 6548 26874
rect 6450 26797 6548 26818
rect 6882 26874 6980 26895
rect 6882 26818 6903 26874
rect 6959 26818 6980 26874
rect 6882 26797 6980 26818
rect 7264 26888 7362 26909
rect 7264 26832 7285 26888
rect 7341 26832 7362 26888
rect 7264 26811 7362 26832
rect 7660 26888 7758 26909
rect 7660 26832 7681 26888
rect 7737 26832 7758 26888
rect 7660 26811 7758 26832
rect 6025 26516 6123 26537
rect 6025 26460 6046 26516
rect 6102 26460 6123 26516
rect 6025 26439 6123 26460
rect 6450 26516 6548 26537
rect 6450 26460 6471 26516
rect 6527 26460 6548 26516
rect 6450 26439 6548 26460
rect 6882 26516 6980 26537
rect 6882 26460 6903 26516
rect 6959 26460 6980 26516
rect 6882 26439 6980 26460
rect 7264 26493 7362 26514
rect 7264 26437 7285 26493
rect 7341 26437 7362 26493
rect 7264 26416 7362 26437
rect 7660 26493 7758 26514
rect 7660 26437 7681 26493
rect 7737 26437 7758 26493
rect 7660 26416 7758 26437
rect 6025 26142 6123 26163
rect 6025 26086 6046 26142
rect 6102 26086 6123 26142
rect 6025 26065 6123 26086
rect 6450 26084 6548 26105
rect 6450 26028 6471 26084
rect 6527 26028 6548 26084
rect 6450 26007 6548 26028
rect 6882 26084 6980 26105
rect 6882 26028 6903 26084
rect 6959 26028 6980 26084
rect 6882 26007 6980 26028
rect 7264 26098 7362 26119
rect 7264 26042 7285 26098
rect 7341 26042 7362 26098
rect 7264 26021 7362 26042
rect 7660 26098 7758 26119
rect 7660 26042 7681 26098
rect 7737 26042 7758 26098
rect 7660 26021 7758 26042
rect 6025 25726 6123 25747
rect 6025 25670 6046 25726
rect 6102 25670 6123 25726
rect 6025 25649 6123 25670
rect 6450 25726 6548 25747
rect 6450 25670 6471 25726
rect 6527 25670 6548 25726
rect 6450 25649 6548 25670
rect 6882 25726 6980 25747
rect 6882 25670 6903 25726
rect 6959 25670 6980 25726
rect 6882 25649 6980 25670
rect 7264 25703 7362 25724
rect 7264 25647 7285 25703
rect 7341 25647 7362 25703
rect 7264 25626 7362 25647
rect 7660 25703 7758 25724
rect 7660 25647 7681 25703
rect 7737 25647 7758 25703
rect 7660 25626 7758 25647
rect 6025 25352 6123 25373
rect 6025 25296 6046 25352
rect 6102 25296 6123 25352
rect 6025 25275 6123 25296
rect 6450 25294 6548 25315
rect 6450 25238 6471 25294
rect 6527 25238 6548 25294
rect 6450 25217 6548 25238
rect 6882 25294 6980 25315
rect 6882 25238 6903 25294
rect 6959 25238 6980 25294
rect 6882 25217 6980 25238
rect 7264 25308 7362 25329
rect 7264 25252 7285 25308
rect 7341 25252 7362 25308
rect 7264 25231 7362 25252
rect 7660 25308 7758 25329
rect 7660 25252 7681 25308
rect 7737 25252 7758 25308
rect 7660 25231 7758 25252
rect 6025 24936 6123 24957
rect 6025 24880 6046 24936
rect 6102 24880 6123 24936
rect 6025 24859 6123 24880
rect 6450 24936 6548 24957
rect 6450 24880 6471 24936
rect 6527 24880 6548 24936
rect 6450 24859 6548 24880
rect 6882 24936 6980 24957
rect 6882 24880 6903 24936
rect 6959 24880 6980 24936
rect 6882 24859 6980 24880
rect 7264 24913 7362 24934
rect 7264 24857 7285 24913
rect 7341 24857 7362 24913
rect 7264 24836 7362 24857
rect 7660 24913 7758 24934
rect 7660 24857 7681 24913
rect 7737 24857 7758 24913
rect 7660 24836 7758 24857
rect 6025 24562 6123 24583
rect 6025 24506 6046 24562
rect 6102 24506 6123 24562
rect 6025 24485 6123 24506
rect 6450 24504 6548 24525
rect 6450 24448 6471 24504
rect 6527 24448 6548 24504
rect 6450 24427 6548 24448
rect 6882 24504 6980 24525
rect 6882 24448 6903 24504
rect 6959 24448 6980 24504
rect 6882 24427 6980 24448
rect 7264 24518 7362 24539
rect 7264 24462 7285 24518
rect 7341 24462 7362 24518
rect 7264 24441 7362 24462
rect 7660 24518 7758 24539
rect 7660 24462 7681 24518
rect 7737 24462 7758 24518
rect 7660 24441 7758 24462
rect 6025 24146 6123 24167
rect 6025 24090 6046 24146
rect 6102 24090 6123 24146
rect 6025 24069 6123 24090
rect 6450 24146 6548 24167
rect 6450 24090 6471 24146
rect 6527 24090 6548 24146
rect 6450 24069 6548 24090
rect 6882 24146 6980 24167
rect 6882 24090 6903 24146
rect 6959 24090 6980 24146
rect 6882 24069 6980 24090
rect 7264 24123 7362 24144
rect 7264 24067 7285 24123
rect 7341 24067 7362 24123
rect 7264 24046 7362 24067
rect 7660 24123 7758 24144
rect 7660 24067 7681 24123
rect 7737 24067 7758 24123
rect 7660 24046 7758 24067
rect 6025 23772 6123 23793
rect 6025 23716 6046 23772
rect 6102 23716 6123 23772
rect 6025 23695 6123 23716
rect 6450 23714 6548 23735
rect 6450 23658 6471 23714
rect 6527 23658 6548 23714
rect 6450 23637 6548 23658
rect 6882 23714 6980 23735
rect 6882 23658 6903 23714
rect 6959 23658 6980 23714
rect 6882 23637 6980 23658
rect 7264 23728 7362 23749
rect 7264 23672 7285 23728
rect 7341 23672 7362 23728
rect 7264 23651 7362 23672
rect 7660 23728 7758 23749
rect 7660 23672 7681 23728
rect 7737 23672 7758 23728
rect 7660 23651 7758 23672
rect 6025 23356 6123 23377
rect 6025 23300 6046 23356
rect 6102 23300 6123 23356
rect 6025 23279 6123 23300
rect 6450 23356 6548 23377
rect 6450 23300 6471 23356
rect 6527 23300 6548 23356
rect 6450 23279 6548 23300
rect 6882 23356 6980 23377
rect 6882 23300 6903 23356
rect 6959 23300 6980 23356
rect 6882 23279 6980 23300
rect 7264 23333 7362 23354
rect 7264 23277 7285 23333
rect 7341 23277 7362 23333
rect 7264 23256 7362 23277
rect 7660 23333 7758 23354
rect 7660 23277 7681 23333
rect 7737 23277 7758 23333
rect 7660 23256 7758 23277
rect 6025 22982 6123 23003
rect 6025 22926 6046 22982
rect 6102 22926 6123 22982
rect 6025 22905 6123 22926
rect 6450 22924 6548 22945
rect 6450 22868 6471 22924
rect 6527 22868 6548 22924
rect 6450 22847 6548 22868
rect 6882 22924 6980 22945
rect 6882 22868 6903 22924
rect 6959 22868 6980 22924
rect 6882 22847 6980 22868
rect 7264 22938 7362 22959
rect 7264 22882 7285 22938
rect 7341 22882 7362 22938
rect 7264 22861 7362 22882
rect 7660 22938 7758 22959
rect 7660 22882 7681 22938
rect 7737 22882 7758 22938
rect 7660 22861 7758 22882
rect 6025 22566 6123 22587
rect 6025 22510 6046 22566
rect 6102 22510 6123 22566
rect 6025 22489 6123 22510
rect 6450 22566 6548 22587
rect 6450 22510 6471 22566
rect 6527 22510 6548 22566
rect 6450 22489 6548 22510
rect 6882 22566 6980 22587
rect 6882 22510 6903 22566
rect 6959 22510 6980 22566
rect 6882 22489 6980 22510
rect 7264 22543 7362 22564
rect 7264 22487 7285 22543
rect 7341 22487 7362 22543
rect 7264 22466 7362 22487
rect 7660 22543 7758 22564
rect 7660 22487 7681 22543
rect 7737 22487 7758 22543
rect 7660 22466 7758 22487
rect 6025 22192 6123 22213
rect 6025 22136 6046 22192
rect 6102 22136 6123 22192
rect 6025 22115 6123 22136
rect 6450 22134 6548 22155
rect 6450 22078 6471 22134
rect 6527 22078 6548 22134
rect 6450 22057 6548 22078
rect 6882 22134 6980 22155
rect 6882 22078 6903 22134
rect 6959 22078 6980 22134
rect 6882 22057 6980 22078
rect 7264 22148 7362 22169
rect 7264 22092 7285 22148
rect 7341 22092 7362 22148
rect 7264 22071 7362 22092
rect 7660 22148 7758 22169
rect 7660 22092 7681 22148
rect 7737 22092 7758 22148
rect 7660 22071 7758 22092
rect 6025 21776 6123 21797
rect 6025 21720 6046 21776
rect 6102 21720 6123 21776
rect 6025 21699 6123 21720
rect 6450 21776 6548 21797
rect 6450 21720 6471 21776
rect 6527 21720 6548 21776
rect 6450 21699 6548 21720
rect 6882 21776 6980 21797
rect 6882 21720 6903 21776
rect 6959 21720 6980 21776
rect 6882 21699 6980 21720
rect 7264 21753 7362 21774
rect 7264 21697 7285 21753
rect 7341 21697 7362 21753
rect 7264 21676 7362 21697
rect 7660 21753 7758 21774
rect 7660 21697 7681 21753
rect 7737 21697 7758 21753
rect 7660 21676 7758 21697
rect 6025 21402 6123 21423
rect 6025 21346 6046 21402
rect 6102 21346 6123 21402
rect 6025 21325 6123 21346
rect 6450 21344 6548 21365
rect 6450 21288 6471 21344
rect 6527 21288 6548 21344
rect 6450 21267 6548 21288
rect 6882 21344 6980 21365
rect 6882 21288 6903 21344
rect 6959 21288 6980 21344
rect 6882 21267 6980 21288
rect 7264 21358 7362 21379
rect 7264 21302 7285 21358
rect 7341 21302 7362 21358
rect 7264 21281 7362 21302
rect 7660 21358 7758 21379
rect 7660 21302 7681 21358
rect 7737 21302 7758 21358
rect 7660 21281 7758 21302
rect 6025 20986 6123 21007
rect 6025 20930 6046 20986
rect 6102 20930 6123 20986
rect 6025 20909 6123 20930
rect 6450 20986 6548 21007
rect 6450 20930 6471 20986
rect 6527 20930 6548 20986
rect 6450 20909 6548 20930
rect 6882 20986 6980 21007
rect 6882 20930 6903 20986
rect 6959 20930 6980 20986
rect 6882 20909 6980 20930
rect 7264 20963 7362 20984
rect 7264 20907 7285 20963
rect 7341 20907 7362 20963
rect 7264 20886 7362 20907
rect 7660 20963 7758 20984
rect 7660 20907 7681 20963
rect 7737 20907 7758 20963
rect 7660 20886 7758 20907
rect 6025 20612 6123 20633
rect 6025 20556 6046 20612
rect 6102 20556 6123 20612
rect 6025 20535 6123 20556
rect 6450 20554 6548 20575
rect 6450 20498 6471 20554
rect 6527 20498 6548 20554
rect 6450 20477 6548 20498
rect 6882 20554 6980 20575
rect 6882 20498 6903 20554
rect 6959 20498 6980 20554
rect 6882 20477 6980 20498
rect 7264 20568 7362 20589
rect 7264 20512 7285 20568
rect 7341 20512 7362 20568
rect 7264 20491 7362 20512
rect 7660 20568 7758 20589
rect 7660 20512 7681 20568
rect 7737 20512 7758 20568
rect 7660 20491 7758 20512
rect 6025 20196 6123 20217
rect 6025 20140 6046 20196
rect 6102 20140 6123 20196
rect 6025 20119 6123 20140
rect 6450 20196 6548 20217
rect 6450 20140 6471 20196
rect 6527 20140 6548 20196
rect 6450 20119 6548 20140
rect 6882 20196 6980 20217
rect 6882 20140 6903 20196
rect 6959 20140 6980 20196
rect 6882 20119 6980 20140
rect 7264 20173 7362 20194
rect 7264 20117 7285 20173
rect 7341 20117 7362 20173
rect 7264 20096 7362 20117
rect 7660 20173 7758 20194
rect 7660 20117 7681 20173
rect 7737 20117 7758 20173
rect 7660 20096 7758 20117
rect 6025 19822 6123 19843
rect 6025 19766 6046 19822
rect 6102 19766 6123 19822
rect 6025 19745 6123 19766
rect 6450 19764 6548 19785
rect 6450 19708 6471 19764
rect 6527 19708 6548 19764
rect 6450 19687 6548 19708
rect 6882 19764 6980 19785
rect 6882 19708 6903 19764
rect 6959 19708 6980 19764
rect 6882 19687 6980 19708
rect 7264 19778 7362 19799
rect 7264 19722 7285 19778
rect 7341 19722 7362 19778
rect 7264 19701 7362 19722
rect 7660 19778 7758 19799
rect 7660 19722 7681 19778
rect 7737 19722 7758 19778
rect 7660 19701 7758 19722
rect 6025 19406 6123 19427
rect 6025 19350 6046 19406
rect 6102 19350 6123 19406
rect 6025 19329 6123 19350
rect 6450 19406 6548 19427
rect 6450 19350 6471 19406
rect 6527 19350 6548 19406
rect 6450 19329 6548 19350
rect 6882 19406 6980 19427
rect 6882 19350 6903 19406
rect 6959 19350 6980 19406
rect 6882 19329 6980 19350
rect 7264 19383 7362 19404
rect 7264 19327 7285 19383
rect 7341 19327 7362 19383
rect 7264 19306 7362 19327
rect 7660 19383 7758 19404
rect 7660 19327 7681 19383
rect 7737 19327 7758 19383
rect 7660 19306 7758 19327
rect 6025 19032 6123 19053
rect 6025 18976 6046 19032
rect 6102 18976 6123 19032
rect 6025 18955 6123 18976
rect 6450 18974 6548 18995
rect 6450 18918 6471 18974
rect 6527 18918 6548 18974
rect 6450 18897 6548 18918
rect 6882 18974 6980 18995
rect 6882 18918 6903 18974
rect 6959 18918 6980 18974
rect 6882 18897 6980 18918
rect 7264 18988 7362 19009
rect 7264 18932 7285 18988
rect 7341 18932 7362 18988
rect 7264 18911 7362 18932
rect 7660 18988 7758 19009
rect 7660 18932 7681 18988
rect 7737 18932 7758 18988
rect 7660 18911 7758 18932
rect 6025 18616 6123 18637
rect 6025 18560 6046 18616
rect 6102 18560 6123 18616
rect 6025 18539 6123 18560
rect 6450 18616 6548 18637
rect 6450 18560 6471 18616
rect 6527 18560 6548 18616
rect 6450 18539 6548 18560
rect 6882 18616 6980 18637
rect 6882 18560 6903 18616
rect 6959 18560 6980 18616
rect 6882 18539 6980 18560
rect 7264 18593 7362 18614
rect 7264 18537 7285 18593
rect 7341 18537 7362 18593
rect 7264 18516 7362 18537
rect 7660 18593 7758 18614
rect 7660 18537 7681 18593
rect 7737 18537 7758 18593
rect 7660 18516 7758 18537
rect 6025 18242 6123 18263
rect 6025 18186 6046 18242
rect 6102 18186 6123 18242
rect 6025 18165 6123 18186
rect 6450 18184 6548 18205
rect 6450 18128 6471 18184
rect 6527 18128 6548 18184
rect 6450 18107 6548 18128
rect 6882 18184 6980 18205
rect 6882 18128 6903 18184
rect 6959 18128 6980 18184
rect 6882 18107 6980 18128
rect 7264 18198 7362 18219
rect 7264 18142 7285 18198
rect 7341 18142 7362 18198
rect 7264 18121 7362 18142
rect 7660 18198 7758 18219
rect 7660 18142 7681 18198
rect 7737 18142 7758 18198
rect 7660 18121 7758 18142
rect 6025 17826 6123 17847
rect 6025 17770 6046 17826
rect 6102 17770 6123 17826
rect 6025 17749 6123 17770
rect 6450 17826 6548 17847
rect 6450 17770 6471 17826
rect 6527 17770 6548 17826
rect 6450 17749 6548 17770
rect 6882 17826 6980 17847
rect 6882 17770 6903 17826
rect 6959 17770 6980 17826
rect 6882 17749 6980 17770
rect 7264 17803 7362 17824
rect 7264 17747 7285 17803
rect 7341 17747 7362 17803
rect 7264 17726 7362 17747
rect 7660 17803 7758 17824
rect 7660 17747 7681 17803
rect 7737 17747 7758 17803
rect 7660 17726 7758 17747
rect 6025 17452 6123 17473
rect 6025 17396 6046 17452
rect 6102 17396 6123 17452
rect 6025 17375 6123 17396
rect 6450 17394 6548 17415
rect 6450 17338 6471 17394
rect 6527 17338 6548 17394
rect 6450 17317 6548 17338
rect 6882 17394 6980 17415
rect 6882 17338 6903 17394
rect 6959 17338 6980 17394
rect 6882 17317 6980 17338
rect 7264 17408 7362 17429
rect 7264 17352 7285 17408
rect 7341 17352 7362 17408
rect 7264 17331 7362 17352
rect 7660 17408 7758 17429
rect 7660 17352 7681 17408
rect 7737 17352 7758 17408
rect 7660 17331 7758 17352
rect 6025 17036 6123 17057
rect 6025 16980 6046 17036
rect 6102 16980 6123 17036
rect 6025 16959 6123 16980
rect 6450 17036 6548 17057
rect 6450 16980 6471 17036
rect 6527 16980 6548 17036
rect 6450 16959 6548 16980
rect 6882 17036 6980 17057
rect 6882 16980 6903 17036
rect 6959 16980 6980 17036
rect 6882 16959 6980 16980
rect 7264 17013 7362 17034
rect 7264 16957 7285 17013
rect 7341 16957 7362 17013
rect 7264 16936 7362 16957
rect 7660 17013 7758 17034
rect 7660 16957 7681 17013
rect 7737 16957 7758 17013
rect 7660 16936 7758 16957
rect 6025 16662 6123 16683
rect 6025 16606 6046 16662
rect 6102 16606 6123 16662
rect 6025 16585 6123 16606
rect 6450 16604 6548 16625
rect 6450 16548 6471 16604
rect 6527 16548 6548 16604
rect 6450 16527 6548 16548
rect 6882 16604 6980 16625
rect 6882 16548 6903 16604
rect 6959 16548 6980 16604
rect 6882 16527 6980 16548
rect 7264 16618 7362 16639
rect 7264 16562 7285 16618
rect 7341 16562 7362 16618
rect 7264 16541 7362 16562
rect 7660 16618 7758 16639
rect 7660 16562 7681 16618
rect 7737 16562 7758 16618
rect 7660 16541 7758 16562
rect 6025 16246 6123 16267
rect 6025 16190 6046 16246
rect 6102 16190 6123 16246
rect 6025 16169 6123 16190
rect 6450 16246 6548 16267
rect 6450 16190 6471 16246
rect 6527 16190 6548 16246
rect 6450 16169 6548 16190
rect 6882 16246 6980 16267
rect 6882 16190 6903 16246
rect 6959 16190 6980 16246
rect 6882 16169 6980 16190
rect 7264 16223 7362 16244
rect 7264 16167 7285 16223
rect 7341 16167 7362 16223
rect 7264 16146 7362 16167
rect 7660 16223 7758 16244
rect 7660 16167 7681 16223
rect 7737 16167 7758 16223
rect 7660 16146 7758 16167
rect 6025 15872 6123 15893
rect 6025 15816 6046 15872
rect 6102 15816 6123 15872
rect 6025 15795 6123 15816
rect 6450 15814 6548 15835
rect 6450 15758 6471 15814
rect 6527 15758 6548 15814
rect 6450 15737 6548 15758
rect 6882 15814 6980 15835
rect 6882 15758 6903 15814
rect 6959 15758 6980 15814
rect 6882 15737 6980 15758
rect 7264 15828 7362 15849
rect 7264 15772 7285 15828
rect 7341 15772 7362 15828
rect 7264 15751 7362 15772
rect 7660 15828 7758 15849
rect 7660 15772 7681 15828
rect 7737 15772 7758 15828
rect 7660 15751 7758 15772
rect 6025 15456 6123 15477
rect 6025 15400 6046 15456
rect 6102 15400 6123 15456
rect 6025 15379 6123 15400
rect 6450 15456 6548 15477
rect 6450 15400 6471 15456
rect 6527 15400 6548 15456
rect 6450 15379 6548 15400
rect 6882 15456 6980 15477
rect 6882 15400 6903 15456
rect 6959 15400 6980 15456
rect 6882 15379 6980 15400
rect 7264 15433 7362 15454
rect 7264 15377 7285 15433
rect 7341 15377 7362 15433
rect 7264 15356 7362 15377
rect 7660 15433 7758 15454
rect 7660 15377 7681 15433
rect 7737 15377 7758 15433
rect 7660 15356 7758 15377
rect 6025 15082 6123 15103
rect 6025 15026 6046 15082
rect 6102 15026 6123 15082
rect 6025 15005 6123 15026
rect 6450 15024 6548 15045
rect 6450 14968 6471 15024
rect 6527 14968 6548 15024
rect 6450 14947 6548 14968
rect 6882 15024 6980 15045
rect 6882 14968 6903 15024
rect 6959 14968 6980 15024
rect 6882 14947 6980 14968
rect 7264 15038 7362 15059
rect 7264 14982 7285 15038
rect 7341 14982 7362 15038
rect 7264 14961 7362 14982
rect 7660 15038 7758 15059
rect 7660 14982 7681 15038
rect 7737 14982 7758 15038
rect 7660 14961 7758 14982
rect 6025 14666 6123 14687
rect 6025 14610 6046 14666
rect 6102 14610 6123 14666
rect 6025 14589 6123 14610
rect 6450 14666 6548 14687
rect 6450 14610 6471 14666
rect 6527 14610 6548 14666
rect 6450 14589 6548 14610
rect 6882 14666 6980 14687
rect 6882 14610 6903 14666
rect 6959 14610 6980 14666
rect 6882 14589 6980 14610
rect 7264 14643 7362 14664
rect 7264 14587 7285 14643
rect 7341 14587 7362 14643
rect 7264 14566 7362 14587
rect 7660 14643 7758 14664
rect 7660 14587 7681 14643
rect 7737 14587 7758 14643
rect 7660 14566 7758 14587
rect 6025 14292 6123 14313
rect 6025 14236 6046 14292
rect 6102 14236 6123 14292
rect 6025 14215 6123 14236
rect 6450 14234 6548 14255
rect 6450 14178 6471 14234
rect 6527 14178 6548 14234
rect 6450 14157 6548 14178
rect 6882 14234 6980 14255
rect 6882 14178 6903 14234
rect 6959 14178 6980 14234
rect 6882 14157 6980 14178
rect 7264 14248 7362 14269
rect 7264 14192 7285 14248
rect 7341 14192 7362 14248
rect 7264 14171 7362 14192
rect 7660 14248 7758 14269
rect 7660 14192 7681 14248
rect 7737 14192 7758 14248
rect 7660 14171 7758 14192
rect 6025 13876 6123 13897
rect 6025 13820 6046 13876
rect 6102 13820 6123 13876
rect 6025 13799 6123 13820
rect 6450 13876 6548 13897
rect 6450 13820 6471 13876
rect 6527 13820 6548 13876
rect 6450 13799 6548 13820
rect 6882 13876 6980 13897
rect 6882 13820 6903 13876
rect 6959 13820 6980 13876
rect 6882 13799 6980 13820
rect 7264 13853 7362 13874
rect 7264 13797 7285 13853
rect 7341 13797 7362 13853
rect 7264 13776 7362 13797
rect 7660 13853 7758 13874
rect 7660 13797 7681 13853
rect 7737 13797 7758 13853
rect 7660 13776 7758 13797
rect 6025 13502 6123 13523
rect 6025 13446 6046 13502
rect 6102 13446 6123 13502
rect 6025 13425 6123 13446
rect 6450 13444 6548 13465
rect 6450 13388 6471 13444
rect 6527 13388 6548 13444
rect 6450 13367 6548 13388
rect 6882 13444 6980 13465
rect 6882 13388 6903 13444
rect 6959 13388 6980 13444
rect 6882 13367 6980 13388
rect 7264 13458 7362 13479
rect 7264 13402 7285 13458
rect 7341 13402 7362 13458
rect 7264 13381 7362 13402
rect 7660 13458 7758 13479
rect 7660 13402 7681 13458
rect 7737 13402 7758 13458
rect 7660 13381 7758 13402
rect 6025 13086 6123 13107
rect 6025 13030 6046 13086
rect 6102 13030 6123 13086
rect 6025 13009 6123 13030
rect 6450 13086 6548 13107
rect 6450 13030 6471 13086
rect 6527 13030 6548 13086
rect 6450 13009 6548 13030
rect 6882 13086 6980 13107
rect 6882 13030 6903 13086
rect 6959 13030 6980 13086
rect 6882 13009 6980 13030
rect 7264 13063 7362 13084
rect 7264 13007 7285 13063
rect 7341 13007 7362 13063
rect 7264 12986 7362 13007
rect 7660 13063 7758 13084
rect 7660 13007 7681 13063
rect 7737 13007 7758 13063
rect 7660 12986 7758 13007
rect 6025 12712 6123 12733
rect 6025 12656 6046 12712
rect 6102 12656 6123 12712
rect 6025 12635 6123 12656
rect 6450 12654 6548 12675
rect 6450 12598 6471 12654
rect 6527 12598 6548 12654
rect 6450 12577 6548 12598
rect 6882 12654 6980 12675
rect 6882 12598 6903 12654
rect 6959 12598 6980 12654
rect 6882 12577 6980 12598
rect 7264 12668 7362 12689
rect 7264 12612 7285 12668
rect 7341 12612 7362 12668
rect 7264 12591 7362 12612
rect 7660 12668 7758 12689
rect 7660 12612 7681 12668
rect 7737 12612 7758 12668
rect 7660 12591 7758 12612
rect 6025 12296 6123 12317
rect 6025 12240 6046 12296
rect 6102 12240 6123 12296
rect 6025 12219 6123 12240
rect 6450 12296 6548 12317
rect 6450 12240 6471 12296
rect 6527 12240 6548 12296
rect 6450 12219 6548 12240
rect 6882 12296 6980 12317
rect 6882 12240 6903 12296
rect 6959 12240 6980 12296
rect 6882 12219 6980 12240
rect 7264 12273 7362 12294
rect 7264 12217 7285 12273
rect 7341 12217 7362 12273
rect 7264 12196 7362 12217
rect 7660 12273 7758 12294
rect 7660 12217 7681 12273
rect 7737 12217 7758 12273
rect 7660 12196 7758 12217
rect 6025 11922 6123 11943
rect 6025 11866 6046 11922
rect 6102 11866 6123 11922
rect 6025 11845 6123 11866
rect 6450 11864 6548 11885
rect 6450 11808 6471 11864
rect 6527 11808 6548 11864
rect 6450 11787 6548 11808
rect 6882 11864 6980 11885
rect 6882 11808 6903 11864
rect 6959 11808 6980 11864
rect 6882 11787 6980 11808
rect 7264 11878 7362 11899
rect 7264 11822 7285 11878
rect 7341 11822 7362 11878
rect 7264 11801 7362 11822
rect 7660 11878 7758 11899
rect 7660 11822 7681 11878
rect 7737 11822 7758 11878
rect 7660 11801 7758 11822
rect 6025 11506 6123 11527
rect 6025 11450 6046 11506
rect 6102 11450 6123 11506
rect 6025 11429 6123 11450
rect 6450 11506 6548 11527
rect 6450 11450 6471 11506
rect 6527 11450 6548 11506
rect 6450 11429 6548 11450
rect 6882 11506 6980 11527
rect 6882 11450 6903 11506
rect 6959 11450 6980 11506
rect 6882 11429 6980 11450
rect 7264 11483 7362 11504
rect 7264 11427 7285 11483
rect 7341 11427 7362 11483
rect 7264 11406 7362 11427
rect 7660 11483 7758 11504
rect 7660 11427 7681 11483
rect 7737 11427 7758 11483
rect 7660 11406 7758 11427
rect 6025 11132 6123 11153
rect 6025 11076 6046 11132
rect 6102 11076 6123 11132
rect 6025 11055 6123 11076
rect 6450 11074 6548 11095
rect 6450 11018 6471 11074
rect 6527 11018 6548 11074
rect 6450 10997 6548 11018
rect 6882 11074 6980 11095
rect 6882 11018 6903 11074
rect 6959 11018 6980 11074
rect 6882 10997 6980 11018
rect 7264 11088 7362 11109
rect 7264 11032 7285 11088
rect 7341 11032 7362 11088
rect 7264 11011 7362 11032
rect 7660 11088 7758 11109
rect 7660 11032 7681 11088
rect 7737 11032 7758 11088
rect 7660 11011 7758 11032
rect 6025 10716 6123 10737
rect 6025 10660 6046 10716
rect 6102 10660 6123 10716
rect 6025 10639 6123 10660
rect 6450 10716 6548 10737
rect 6450 10660 6471 10716
rect 6527 10660 6548 10716
rect 6450 10639 6548 10660
rect 6882 10716 6980 10737
rect 6882 10660 6903 10716
rect 6959 10660 6980 10716
rect 6882 10639 6980 10660
rect 7264 10693 7362 10714
rect 7264 10637 7285 10693
rect 7341 10637 7362 10693
rect 7264 10616 7362 10637
rect 7660 10693 7758 10714
rect 7660 10637 7681 10693
rect 7737 10637 7758 10693
rect 7660 10616 7758 10637
rect 6025 10342 6123 10363
rect 6025 10286 6046 10342
rect 6102 10286 6123 10342
rect 6025 10265 6123 10286
rect 6450 10284 6548 10305
rect 6450 10228 6471 10284
rect 6527 10228 6548 10284
rect 6450 10207 6548 10228
rect 6882 10284 6980 10305
rect 6882 10228 6903 10284
rect 6959 10228 6980 10284
rect 6882 10207 6980 10228
rect 7264 10298 7362 10319
rect 7264 10242 7285 10298
rect 7341 10242 7362 10298
rect 7264 10221 7362 10242
rect 7660 10298 7758 10319
rect 7660 10242 7681 10298
rect 7737 10242 7758 10298
rect 7660 10221 7758 10242
rect 6025 9926 6123 9947
rect 6025 9870 6046 9926
rect 6102 9870 6123 9926
rect 6025 9849 6123 9870
rect 6450 9926 6548 9947
rect 6450 9870 6471 9926
rect 6527 9870 6548 9926
rect 6450 9849 6548 9870
rect 6882 9926 6980 9947
rect 6882 9870 6903 9926
rect 6959 9870 6980 9926
rect 6882 9849 6980 9870
rect 7264 9903 7362 9924
rect 7264 9847 7285 9903
rect 7341 9847 7362 9903
rect 7264 9826 7362 9847
rect 7660 9903 7758 9924
rect 7660 9847 7681 9903
rect 7737 9847 7758 9903
rect 7660 9826 7758 9847
rect 6025 9552 6123 9573
rect 6025 9496 6046 9552
rect 6102 9496 6123 9552
rect 6025 9475 6123 9496
rect 6450 9494 6548 9515
rect 6450 9438 6471 9494
rect 6527 9438 6548 9494
rect 6450 9417 6548 9438
rect 6882 9494 6980 9515
rect 6882 9438 6903 9494
rect 6959 9438 6980 9494
rect 6882 9417 6980 9438
rect 7264 9508 7362 9529
rect 7264 9452 7285 9508
rect 7341 9452 7362 9508
rect 7264 9431 7362 9452
rect 7660 9508 7758 9529
rect 7660 9452 7681 9508
rect 7737 9452 7758 9508
rect 7660 9431 7758 9452
rect 6025 9136 6123 9157
rect 6025 9080 6046 9136
rect 6102 9080 6123 9136
rect 6025 9059 6123 9080
rect 6450 9136 6548 9157
rect 6450 9080 6471 9136
rect 6527 9080 6548 9136
rect 6450 9059 6548 9080
rect 6882 9136 6980 9157
rect 6882 9080 6903 9136
rect 6959 9080 6980 9136
rect 6882 9059 6980 9080
rect 7264 9113 7362 9134
rect 7264 9057 7285 9113
rect 7341 9057 7362 9113
rect 7264 9036 7362 9057
rect 7660 9113 7758 9134
rect 7660 9057 7681 9113
rect 7737 9057 7758 9113
rect 7660 9036 7758 9057
rect 6025 8762 6123 8783
rect 6025 8706 6046 8762
rect 6102 8706 6123 8762
rect 6025 8685 6123 8706
rect 6450 8704 6548 8725
rect 6450 8648 6471 8704
rect 6527 8648 6548 8704
rect 6450 8627 6548 8648
rect 6882 8704 6980 8725
rect 6882 8648 6903 8704
rect 6959 8648 6980 8704
rect 6882 8627 6980 8648
rect 7264 8718 7362 8739
rect 7264 8662 7285 8718
rect 7341 8662 7362 8718
rect 7264 8641 7362 8662
rect 7660 8718 7758 8739
rect 7660 8662 7681 8718
rect 7737 8662 7758 8718
rect 7660 8641 7758 8662
rect 6025 8346 6123 8367
rect 6025 8290 6046 8346
rect 6102 8290 6123 8346
rect 6025 8269 6123 8290
rect 6450 8346 6548 8367
rect 6450 8290 6471 8346
rect 6527 8290 6548 8346
rect 6450 8269 6548 8290
rect 6882 8346 6980 8367
rect 6882 8290 6903 8346
rect 6959 8290 6980 8346
rect 6882 8269 6980 8290
rect 7264 8323 7362 8344
rect 7264 8267 7285 8323
rect 7341 8267 7362 8323
rect 7264 8246 7362 8267
rect 7660 8323 7758 8344
rect 7660 8267 7681 8323
rect 7737 8267 7758 8323
rect 7660 8246 7758 8267
rect 6025 7972 6123 7993
rect 6025 7916 6046 7972
rect 6102 7916 6123 7972
rect 6025 7895 6123 7916
rect 6450 7914 6548 7935
rect 6450 7858 6471 7914
rect 6527 7858 6548 7914
rect 6450 7837 6548 7858
rect 6882 7914 6980 7935
rect 6882 7858 6903 7914
rect 6959 7858 6980 7914
rect 6882 7837 6980 7858
rect 7264 7928 7362 7949
rect 7264 7872 7285 7928
rect 7341 7872 7362 7928
rect 7264 7851 7362 7872
rect 7660 7928 7758 7949
rect 7660 7872 7681 7928
rect 7737 7872 7758 7928
rect 7660 7851 7758 7872
rect 2611 7479 2709 7577
rect 3036 7479 3134 7577
rect 3468 7479 3566 7577
rect 6025 7556 6123 7577
rect 3850 7456 3948 7554
rect 4246 7456 4344 7554
rect 6025 7500 6046 7556
rect 6102 7500 6123 7556
rect 6025 7479 6123 7500
rect 6450 7556 6548 7577
rect 6450 7500 6471 7556
rect 6527 7500 6548 7556
rect 6450 7479 6548 7500
rect 6882 7556 6980 7577
rect 6882 7500 6903 7556
rect 6959 7500 6980 7556
rect 6882 7479 6980 7500
rect 7264 7533 7362 7554
rect 7264 7477 7285 7533
rect 7341 7477 7362 7533
rect 7264 7456 7362 7477
rect 7660 7533 7758 7554
rect 7660 7477 7681 7533
rect 7737 7477 7758 7533
rect 7660 7456 7758 7477
rect 6025 7182 6123 7203
rect 6025 7126 6046 7182
rect 6102 7126 6123 7182
rect 6025 7105 6123 7126
rect 6450 7124 6548 7145
rect 6450 7068 6471 7124
rect 6527 7068 6548 7124
rect 6450 7047 6548 7068
rect 6882 7124 6980 7145
rect 6882 7068 6903 7124
rect 6959 7068 6980 7124
rect 6882 7047 6980 7068
rect 7264 7138 7362 7159
rect 7264 7082 7285 7138
rect 7341 7082 7362 7138
rect 7264 7061 7362 7082
rect 7660 7138 7758 7159
rect 7660 7082 7681 7138
rect 7737 7082 7758 7138
rect 7660 7061 7758 7082
rect 2611 6689 2709 6787
rect 3036 6689 3134 6787
rect 3468 6689 3566 6787
rect 6025 6766 6123 6787
rect 3850 6666 3948 6764
rect 4246 6666 4344 6764
rect 6025 6710 6046 6766
rect 6102 6710 6123 6766
rect 6025 6689 6123 6710
rect 6450 6766 6548 6787
rect 6450 6710 6471 6766
rect 6527 6710 6548 6766
rect 6450 6689 6548 6710
rect 6882 6766 6980 6787
rect 6882 6710 6903 6766
rect 6959 6710 6980 6766
rect 6882 6689 6980 6710
rect 7264 6743 7362 6764
rect 7264 6687 7285 6743
rect 7341 6687 7362 6743
rect 7264 6666 7362 6687
rect 7660 6743 7758 6764
rect 7660 6687 7681 6743
rect 7737 6687 7758 6743
rect 7660 6666 7758 6687
rect 6025 6392 6123 6413
rect 6025 6336 6046 6392
rect 6102 6336 6123 6392
rect 6025 6315 6123 6336
rect 6450 6334 6548 6355
rect 6450 6278 6471 6334
rect 6527 6278 6548 6334
rect 6450 6257 6548 6278
rect 6882 6334 6980 6355
rect 6882 6278 6903 6334
rect 6959 6278 6980 6334
rect 6882 6257 6980 6278
rect 7264 6348 7362 6369
rect 7264 6292 7285 6348
rect 7341 6292 7362 6348
rect 7264 6271 7362 6292
rect 7660 6348 7758 6369
rect 7660 6292 7681 6348
rect 7737 6292 7758 6348
rect 7660 6271 7758 6292
rect 2611 5899 2709 5997
rect 3036 5899 3134 5997
rect 3468 5899 3566 5997
rect 6025 5976 6123 5997
rect 3850 5876 3948 5974
rect 4246 5876 4344 5974
rect 6025 5920 6046 5976
rect 6102 5920 6123 5976
rect 6025 5899 6123 5920
rect 6450 5976 6548 5997
rect 6450 5920 6471 5976
rect 6527 5920 6548 5976
rect 6450 5899 6548 5920
rect 6882 5976 6980 5997
rect 6882 5920 6903 5976
rect 6959 5920 6980 5976
rect 6882 5899 6980 5920
rect 7264 5953 7362 5974
rect 7264 5897 7285 5953
rect 7341 5897 7362 5953
rect 7264 5876 7362 5897
rect 7660 5953 7758 5974
rect 7660 5897 7681 5953
rect 7737 5897 7758 5953
rect 7660 5876 7758 5897
rect 6025 5602 6123 5623
rect 6025 5546 6046 5602
rect 6102 5546 6123 5602
rect 6025 5525 6123 5546
rect 6450 5544 6548 5565
rect 6450 5488 6471 5544
rect 6527 5488 6548 5544
rect 6450 5467 6548 5488
rect 6882 5544 6980 5565
rect 6882 5488 6903 5544
rect 6959 5488 6980 5544
rect 6882 5467 6980 5488
rect 7264 5558 7362 5579
rect 7264 5502 7285 5558
rect 7341 5502 7362 5558
rect 7264 5481 7362 5502
rect 7660 5558 7758 5579
rect 7660 5502 7681 5558
rect 7737 5502 7758 5558
rect 7660 5481 7758 5502
rect 1156 5086 1254 5184
rect 1552 5086 1650 5184
rect 2611 5109 2709 5207
rect 3036 5109 3134 5207
rect 3468 5109 3566 5207
rect 6025 5186 6123 5207
rect 3850 5086 3948 5184
rect 4246 5086 4344 5184
rect 6025 5130 6046 5186
rect 6102 5130 6123 5186
rect 6025 5109 6123 5130
rect 6450 5186 6548 5207
rect 6450 5130 6471 5186
rect 6527 5130 6548 5186
rect 6450 5109 6548 5130
rect 6882 5186 6980 5207
rect 6882 5130 6903 5186
rect 6959 5130 6980 5186
rect 6882 5109 6980 5130
rect 7264 5163 7362 5184
rect 7264 5107 7285 5163
rect 7341 5107 7362 5163
rect 7264 5086 7362 5107
rect 7660 5163 7758 5184
rect 7660 5107 7681 5163
rect 7737 5107 7758 5163
rect 7660 5086 7758 5107
rect 6025 4812 6123 4833
rect 6025 4756 6046 4812
rect 6102 4756 6123 4812
rect 6025 4735 6123 4756
rect 6450 4754 6548 4775
rect 6450 4698 6471 4754
rect 6527 4698 6548 4754
rect 6450 4677 6548 4698
rect 6882 4754 6980 4775
rect 6882 4698 6903 4754
rect 6959 4698 6980 4754
rect 6882 4677 6980 4698
rect 7264 4768 7362 4789
rect 7264 4712 7285 4768
rect 7341 4712 7362 4768
rect 7264 4691 7362 4712
rect 7660 4768 7758 4789
rect 7660 4712 7681 4768
rect 7737 4712 7758 4768
rect 7660 4691 7758 4712
rect 6025 4396 6123 4417
rect 6025 4340 6046 4396
rect 6102 4340 6123 4396
rect 6025 4319 6123 4340
rect 6450 4396 6548 4417
rect 6450 4340 6471 4396
rect 6527 4340 6548 4396
rect 6450 4319 6548 4340
rect 6882 4396 6980 4417
rect 6882 4340 6903 4396
rect 6959 4340 6980 4396
rect 6882 4319 6980 4340
rect 7264 4373 7362 4394
rect 7264 4317 7285 4373
rect 7341 4317 7362 4373
rect 7264 4296 7362 4317
rect 7660 4373 7758 4394
rect 7660 4317 7681 4373
rect 7737 4317 7758 4373
rect 7660 4296 7758 4317
rect 6025 4022 6123 4043
rect 6025 3966 6046 4022
rect 6102 3966 6123 4022
rect 6025 3945 6123 3966
rect 6450 3964 6548 3985
rect 6450 3908 6471 3964
rect 6527 3908 6548 3964
rect 6450 3887 6548 3908
rect 6882 3964 6980 3985
rect 6882 3908 6903 3964
rect 6959 3908 6980 3964
rect 6882 3887 6980 3908
rect 7264 3978 7362 3999
rect 7264 3922 7285 3978
rect 7341 3922 7362 3978
rect 7264 3901 7362 3922
rect 7660 3978 7758 3999
rect 7660 3922 7681 3978
rect 7737 3922 7758 3978
rect 7660 3901 7758 3922
rect 3046 3513 3144 3611
rect 3471 3513 3569 3611
rect 6025 3606 6123 3627
rect 3850 3506 3948 3604
rect 4246 3506 4344 3604
rect 6025 3550 6046 3606
rect 6102 3550 6123 3606
rect 6025 3529 6123 3550
rect 6450 3606 6548 3627
rect 6450 3550 6471 3606
rect 6527 3550 6548 3606
rect 6450 3529 6548 3550
rect 6882 3606 6980 3627
rect 6882 3550 6903 3606
rect 6959 3550 6980 3606
rect 6882 3529 6980 3550
rect 7264 3583 7362 3604
rect 7264 3527 7285 3583
rect 7341 3527 7362 3583
rect 7264 3506 7362 3527
rect 7660 3583 7758 3604
rect 7660 3527 7681 3583
rect 7737 3527 7758 3583
rect 7660 3506 7758 3527
rect 6025 3232 6123 3253
rect 6025 3176 6046 3232
rect 6102 3176 6123 3232
rect 6025 3155 6123 3176
rect 6450 3174 6548 3195
rect 6450 3118 6471 3174
rect 6527 3118 6548 3174
rect 6450 3097 6548 3118
rect 6882 3174 6980 3195
rect 6882 3118 6903 3174
rect 6959 3118 6980 3174
rect 6882 3097 6980 3118
rect 7264 3188 7362 3209
rect 7264 3132 7285 3188
rect 7341 3132 7362 3188
rect 7264 3111 7362 3132
rect 7660 3188 7758 3209
rect 7660 3132 7681 3188
rect 7737 3132 7758 3188
rect 7660 3111 7758 3132
rect 1752 2716 1850 2814
rect 2148 2716 2246 2814
rect 3046 2723 3144 2821
rect 3471 2723 3569 2821
rect 6025 2816 6123 2837
rect 3850 2716 3948 2814
rect 4246 2716 4344 2814
rect 6025 2760 6046 2816
rect 6102 2760 6123 2816
rect 6025 2739 6123 2760
rect 6450 2816 6548 2837
rect 6450 2760 6471 2816
rect 6527 2760 6548 2816
rect 6450 2739 6548 2760
rect 6882 2816 6980 2837
rect 6882 2760 6903 2816
rect 6959 2760 6980 2816
rect 6882 2739 6980 2760
rect 7264 2793 7362 2814
rect 7264 2737 7285 2793
rect 7341 2737 7362 2793
rect 7264 2716 7362 2737
rect 7660 2793 7758 2814
rect 7660 2737 7681 2793
rect 7737 2737 7758 2793
rect 7660 2716 7758 2737
rect 6025 2442 6123 2463
rect 6025 2386 6046 2442
rect 6102 2386 6123 2442
rect 6025 2365 6123 2386
rect 6450 2384 6548 2405
rect 6450 2328 6471 2384
rect 6527 2328 6548 2384
rect 6450 2307 6548 2328
rect 6882 2384 6980 2405
rect 6882 2328 6903 2384
rect 6959 2328 6980 2384
rect 6882 2307 6980 2328
rect 7264 2398 7362 2419
rect 7264 2342 7285 2398
rect 7341 2342 7362 2398
rect 7264 2321 7362 2342
rect 7660 2398 7758 2419
rect 7660 2342 7681 2398
rect 7737 2342 7758 2398
rect 7660 2321 7758 2342
rect 6025 2026 6123 2047
rect 6025 1970 6046 2026
rect 6102 1970 6123 2026
rect 6025 1949 6123 1970
rect 6450 2026 6548 2047
rect 6450 1970 6471 2026
rect 6527 1970 6548 2026
rect 6450 1949 6548 1970
rect 6882 2026 6980 2047
rect 6882 1970 6903 2026
rect 6959 1970 6980 2026
rect 6882 1949 6980 1970
rect 7264 2003 7362 2024
rect 7264 1947 7285 2003
rect 7341 1947 7362 2003
rect 7264 1926 7362 1947
rect 7660 2003 7758 2024
rect 7660 1947 7681 2003
rect 7737 1947 7758 2003
rect 7660 1926 7758 1947
rect 6025 1652 6123 1673
rect 6025 1596 6046 1652
rect 6102 1596 6123 1652
rect 6025 1575 6123 1596
rect 6450 1594 6548 1615
rect 6450 1538 6471 1594
rect 6527 1538 6548 1594
rect 6450 1517 6548 1538
rect 6882 1594 6980 1615
rect 6882 1538 6903 1594
rect 6959 1538 6980 1594
rect 6882 1517 6980 1538
rect 7264 1608 7362 1629
rect 7264 1552 7285 1608
rect 7341 1552 7362 1608
rect 7264 1531 7362 1552
rect 7660 1608 7758 1629
rect 7660 1552 7681 1608
rect 7737 1552 7758 1608
rect 7660 1531 7758 1552
rect 3046 1143 3144 1241
rect 3471 1143 3569 1241
rect 6025 1236 6123 1257
rect 3850 1136 3948 1234
rect 4246 1136 4344 1234
rect 6025 1180 6046 1236
rect 6102 1180 6123 1236
rect 6025 1159 6123 1180
rect 6450 1236 6548 1257
rect 6450 1180 6471 1236
rect 6527 1180 6548 1236
rect 6450 1159 6548 1180
rect 6882 1236 6980 1257
rect 6882 1180 6903 1236
rect 6959 1180 6980 1236
rect 6882 1159 6980 1180
rect 7264 1213 7362 1234
rect 7264 1157 7285 1213
rect 7341 1157 7362 1213
rect 7264 1136 7362 1157
rect 7660 1213 7758 1234
rect 7660 1157 7681 1213
rect 7737 1157 7758 1213
rect 7660 1136 7758 1157
rect 6025 862 6123 883
rect 6025 806 6046 862
rect 6102 806 6123 862
rect 6025 785 6123 806
rect 6450 804 6548 825
rect 6450 748 6471 804
rect 6527 748 6548 804
rect 6450 727 6548 748
rect 6882 804 6980 825
rect 6882 748 6903 804
rect 6959 748 6980 804
rect 6882 727 6980 748
rect 7264 818 7362 839
rect 7264 762 7285 818
rect 7341 762 7362 818
rect 7264 741 7362 762
rect 7660 818 7758 839
rect 7660 762 7681 818
rect 7737 762 7758 818
rect 7660 741 7758 762
rect 1752 346 1850 444
rect 2148 346 2246 444
rect 3046 353 3144 451
rect 3471 353 3569 451
rect 6025 446 6123 467
rect 3850 346 3948 444
rect 4246 346 4344 444
rect 6025 390 6046 446
rect 6102 390 6123 446
rect 6025 369 6123 390
rect 6450 446 6548 467
rect 6450 390 6471 446
rect 6527 390 6548 446
rect 6450 369 6548 390
rect 6882 446 6980 467
rect 6882 390 6903 446
rect 6959 390 6980 446
rect 6882 369 6980 390
rect 7264 423 7362 444
rect 7264 367 7285 423
rect 7341 367 7362 423
rect 7264 346 7362 367
rect 7660 423 7758 444
rect 7660 367 7681 423
rect 7737 367 7758 423
rect 7660 346 7758 367
use contact_17  contact_17_389
timestamp 1624857261
transform 1 0 80 0 1 591
box 0 0 1 1
use contact_14  contact_14_21
timestamp 1624857261
transform 1 0 1428 0 1 587
box 0 0 1 1
use contact_17  contact_17_390
timestamp 1624857261
transform 1 0 0 0 1 141
box 0 0 1 1
use contact_14  contact_14_22
timestamp 1624857261
transform 1 0 1348 0 1 137
box 0 0 1 1
use contact_17  contact_17_387
timestamp 1624857261
transform 1 0 240 0 1 2961
box 0 0 1 1
use contact_14  contact_14_19
timestamp 1624857261
transform 1 0 1428 0 1 2957
box 0 0 1 1
use contact_17  contact_17_388
timestamp 1624857261
transform 1 0 160 0 1 2511
box 0 0 1 1
use contact_14  contact_14_20
timestamp 1624857261
transform 1 0 1348 0 1 2507
box 0 0 1 1
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1624857261
transform 1 0 1283 0 1 2370
box 61 -56 3178 1636
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1624857261
transform 1 0 1283 0 1 0
box 61 -56 3178 1636
use contact_14  contact_14_15
timestamp 1624857261
transform 1 0 4414 0 1 87
box 0 0 1 1
use contact_19  contact_19_650
timestamp 1624857261
transform 1 0 4411 0 1 88
box 0 0 1 1
use contact_20  contact_20_15
timestamp 1624857261
transform 1 0 4505 0 1 -32
box 0 0 1 1
use contact_17  contact_17_383
timestamp 1624857261
transform 1 0 4504 0 1 52
box 0 0 1 1
use contact_17  contact_17_382
timestamp 1624857261
transform 1 0 4824 0 1 164
box 0 0 1 1
use contact_20  contact_20_14
timestamp 1624857261
transform 1 0 4585 0 1 363
box 0 0 1 1
use contact_17  contact_17_378
timestamp 1624857261
transform 1 0 5144 0 1 478
box 0 0 1 1
use contact_17  contact_17_381
timestamp 1624857261
transform 1 0 5144 0 1 254
box 0 0 1 1
use contact_7  contact_7_253
timestamp 1624857261
transform 1 0 6041 0 1 381
box 0 0 1 1
use contact_19  contact_19_253
timestamp 1624857261
transform 1 0 6042 0 1 386
box 0 0 1 1
use contact_7  contact_7_634
timestamp 1624857261
transform 1 0 6466 0 1 381
box 0 0 1 1
use contact_19  contact_19_634
timestamp 1624857261
transform 1 0 6467 0 1 386
box 0 0 1 1
use contact_7  contact_7_632
timestamp 1624857261
transform 1 0 6898 0 1 381
box 0 0 1 1
use contact_19  contact_19_632
timestamp 1624857261
transform 1 0 6899 0 1 386
box 0 0 1 1
use contact_7  contact_7_252
timestamp 1624857261
transform 1 0 7280 0 1 358
box 0 0 1 1
use contact_19  contact_19_252
timestamp 1624857261
transform 1 0 7281 0 1 363
box 0 0 1 1
use and3_dec  and3_dec_127
timestamp 1624857261
transform 1 0 5803 0 1 0
box 0 -60 2072 490
use and3_dec  and3_dec_126
timestamp 1624857261
transform 1 0 5803 0 -1 790
box 0 -60 2072 490
use contact_19  contact_19_649
timestamp 1624857261
transform 1 0 4411 0 1 638
box 0 0 1 1
use contact_14  contact_14_14
timestamp 1624857261
transform 1 0 4414 0 1 637
box 0 0 1 1
use contact_17  contact_17_379
timestamp 1624857261
transform 1 0 4824 0 1 568
box 0 0 1 1
use contact_17  contact_17_380
timestamp 1624857261
transform 1 0 4584 0 1 680
box 0 0 1 1
use contact_20  contact_20_13
timestamp 1624857261
transform 1 0 4665 0 1 758
box 0 0 1 1
use contact_7  contact_7_631
timestamp 1624857261
transform 1 0 6466 0 1 739
box 0 0 1 1
use contact_19  contact_19_631
timestamp 1624857261
transform 1 0 6467 0 1 744
box 0 0 1 1
use contact_7  contact_7_629
timestamp 1624857261
transform 1 0 6898 0 1 739
box 0 0 1 1
use contact_19  contact_19_629
timestamp 1624857261
transform 1 0 6899 0 1 744
box 0 0 1 1
use contact_7  contact_7_250
timestamp 1624857261
transform 1 0 7280 0 1 753
box 0 0 1 1
use contact_19  contact_19_250
timestamp 1624857261
transform 1 0 7281 0 1 758
box 0 0 1 1
use contact_14  contact_14_13
timestamp 1624857261
transform 1 0 4414 0 1 877
box 0 0 1 1
use contact_19  contact_19_648
timestamp 1624857261
transform 1 0 4411 0 1 878
box 0 0 1 1
use contact_17  contact_17_377
timestamp 1624857261
transform 1 0 4664 0 1 842
box 0 0 1 1
use contact_17  contact_17_376
timestamp 1624857261
transform 1 0 4824 0 1 954
box 0 0 1 1
use contact_19  contact_19_251
timestamp 1624857261
transform 1 0 6042 0 1 802
box 0 0 1 1
use contact_7  contact_7_251
timestamp 1624857261
transform 1 0 6041 0 1 797
box 0 0 1 1
use and3_dec  and3_dec_125
timestamp 1624857261
transform 1 0 5803 0 1 790
box 0 -60 2072 490
use contact_20  contact_20_12
timestamp 1624857261
transform 1 0 4745 0 1 1153
box 0 0 1 1
use contact_17  contact_17_372
timestamp 1624857261
transform 1 0 5144 0 1 1268
box 0 0 1 1
use contact_17  contact_17_375
timestamp 1624857261
transform 1 0 5144 0 1 1044
box 0 0 1 1
use contact_7  contact_7_249
timestamp 1624857261
transform 1 0 6041 0 1 1171
box 0 0 1 1
use contact_19  contact_19_249
timestamp 1624857261
transform 1 0 6042 0 1 1176
box 0 0 1 1
use contact_7  contact_7_628
timestamp 1624857261
transform 1 0 6466 0 1 1171
box 0 0 1 1
use contact_19  contact_19_628
timestamp 1624857261
transform 1 0 6467 0 1 1176
box 0 0 1 1
use contact_7  contact_7_626
timestamp 1624857261
transform 1 0 6898 0 1 1171
box 0 0 1 1
use contact_19  contact_19_626
timestamp 1624857261
transform 1 0 6899 0 1 1176
box 0 0 1 1
use contact_7  contact_7_248
timestamp 1624857261
transform 1 0 7280 0 1 1148
box 0 0 1 1
use contact_19  contact_19_248
timestamp 1624857261
transform 1 0 7281 0 1 1153
box 0 0 1 1
use contact_19  contact_19_647
timestamp 1624857261
transform 1 0 4411 0 1 1428
box 0 0 1 1
use contact_14  contact_14_12
timestamp 1624857261
transform 1 0 4414 0 1 1427
box 0 0 1 1
use contact_17  contact_17_373
timestamp 1624857261
transform 1 0 4824 0 1 1358
box 0 0 1 1
use contact_17  contact_17_374
timestamp 1624857261
transform 1 0 4744 0 1 1470
box 0 0 1 1
use contact_7  contact_7_247
timestamp 1624857261
transform 1 0 6041 0 1 1587
box 0 0 1 1
use contact_19  contact_19_247
timestamp 1624857261
transform 1 0 6042 0 1 1592
box 0 0 1 1
use contact_7  contact_7_625
timestamp 1624857261
transform 1 0 6466 0 1 1529
box 0 0 1 1
use contact_19  contact_19_625
timestamp 1624857261
transform 1 0 6467 0 1 1534
box 0 0 1 1
use contact_7  contact_7_623
timestamp 1624857261
transform 1 0 6898 0 1 1529
box 0 0 1 1
use contact_19  contact_19_623
timestamp 1624857261
transform 1 0 6899 0 1 1534
box 0 0 1 1
use contact_7  contact_7_246
timestamp 1624857261
transform 1 0 7280 0 1 1543
box 0 0 1 1
use contact_19  contact_19_246
timestamp 1624857261
transform 1 0 7281 0 1 1548
box 0 0 1 1
use and3_dec  and3_dec_124
timestamp 1624857261
transform 1 0 5803 0 -1 1580
box 0 -60 2072 490
use and3_dec  and3_dec_123
timestamp 1624857261
transform 1 0 5803 0 1 1580
box 0 -60 2072 490
use contact_17  contact_17_371
timestamp 1624857261
transform 1 0 4504 0 1 1632
box 0 0 1 1
use contact_17  contact_17_370
timestamp 1624857261
transform 1 0 4904 0 1 1744
box 0 0 1 1
use contact_17  contact_17_369
timestamp 1624857261
transform 1 0 5144 0 1 1834
box 0 0 1 1
use contact_17  contact_17_366
timestamp 1624857261
transform 1 0 5144 0 1 2058
box 0 0 1 1
use contact_19  contact_19_622
timestamp 1624857261
transform 1 0 6467 0 1 1966
box 0 0 1 1
use contact_7  contact_7_622
timestamp 1624857261
transform 1 0 6466 0 1 1961
box 0 0 1 1
use contact_19  contact_19_620
timestamp 1624857261
transform 1 0 6899 0 1 1966
box 0 0 1 1
use contact_7  contact_7_620
timestamp 1624857261
transform 1 0 6898 0 1 1961
box 0 0 1 1
use contact_19  contact_19_245
timestamp 1624857261
transform 1 0 6042 0 1 1966
box 0 0 1 1
use contact_7  contact_7_245
timestamp 1624857261
transform 1 0 6041 0 1 1961
box 0 0 1 1
use contact_19  contact_19_244
timestamp 1624857261
transform 1 0 7281 0 1 1943
box 0 0 1 1
use contact_7  contact_7_244
timestamp 1624857261
transform 1 0 7280 0 1 1938
box 0 0 1 1
use and3_dec  and3_dec_122
timestamp 1624857261
transform 1 0 5803 0 -1 2370
box 0 -60 2072 490
use contact_17  contact_17_368
timestamp 1624857261
transform 1 0 4584 0 1 2260
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1624857261
transform 1 0 4825 0 1 2338
box 0 0 1 1
use contact_17  contact_17_367
timestamp 1624857261
transform 1 0 4904 0 1 2148
box 0 0 1 1
use contact_7  contact_7_243
timestamp 1624857261
transform 1 0 6041 0 1 2377
box 0 0 1 1
use contact_19  contact_19_243
timestamp 1624857261
transform 1 0 6042 0 1 2382
box 0 0 1 1
use contact_7  contact_7_619
timestamp 1624857261
transform 1 0 6466 0 1 2319
box 0 0 1 1
use contact_19  contact_19_619
timestamp 1624857261
transform 1 0 6467 0 1 2324
box 0 0 1 1
use contact_7  contact_7_617
timestamp 1624857261
transform 1 0 6898 0 1 2319
box 0 0 1 1
use contact_19  contact_19_617
timestamp 1624857261
transform 1 0 6899 0 1 2324
box 0 0 1 1
use contact_7  contact_7_242
timestamp 1624857261
transform 1 0 7280 0 1 2333
box 0 0 1 1
use contact_19  contact_19_242
timestamp 1624857261
transform 1 0 7281 0 1 2338
box 0 0 1 1
use contact_14  contact_14_11
timestamp 1624857261
transform 1 0 4414 0 1 2457
box 0 0 1 1
use contact_19  contact_19_646
timestamp 1624857261
transform 1 0 4411 0 1 2458
box 0 0 1 1
use contact_17  contact_17_365
timestamp 1624857261
transform 1 0 4664 0 1 2422
box 0 0 1 1
use contact_17  contact_17_364
timestamp 1624857261
transform 1 0 4904 0 1 2534
box 0 0 1 1
use contact_17  contact_17_363
timestamp 1624857261
transform 1 0 5144 0 1 2624
box 0 0 1 1
use and3_dec  and3_dec_121
timestamp 1624857261
transform 1 0 5803 0 1 2370
box 0 -60 2072 490
use and3_dec  and3_dec_120
timestamp 1624857261
transform 1 0 5803 0 -1 3160
box 0 -60 2072 490
use contact_17  contact_17_360
timestamp 1624857261
transform 1 0 5144 0 1 2848
box 0 0 1 1
use contact_17  contact_17_361
timestamp 1624857261
transform 1 0 4904 0 1 2938
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1624857261
transform 1 0 4905 0 1 2733
box 0 0 1 1
use contact_7  contact_7_241
timestamp 1624857261
transform 1 0 6041 0 1 2751
box 0 0 1 1
use contact_19  contact_19_241
timestamp 1624857261
transform 1 0 6042 0 1 2756
box 0 0 1 1
use contact_7  contact_7_616
timestamp 1624857261
transform 1 0 6466 0 1 2751
box 0 0 1 1
use contact_19  contact_19_616
timestamp 1624857261
transform 1 0 6467 0 1 2756
box 0 0 1 1
use contact_7  contact_7_614
timestamp 1624857261
transform 1 0 6898 0 1 2751
box 0 0 1 1
use contact_19  contact_19_614
timestamp 1624857261
transform 1 0 6899 0 1 2756
box 0 0 1 1
use contact_7  contact_7_240
timestamp 1624857261
transform 1 0 7280 0 1 2728
box 0 0 1 1
use contact_19  contact_19_240
timestamp 1624857261
transform 1 0 7281 0 1 2733
box 0 0 1 1
use contact_17  contact_17_359
timestamp 1624857261
transform 1 0 4504 0 1 3212
box 0 0 1 1
use contact_19  contact_19_645
timestamp 1624857261
transform 1 0 4411 0 1 3008
box 0 0 1 1
use contact_14  contact_14_10
timestamp 1624857261
transform 1 0 4414 0 1 3007
box 0 0 1 1
use contact_17  contact_17_362
timestamp 1624857261
transform 1 0 4744 0 1 3050
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1624857261
transform 1 0 4985 0 1 3128
box 0 0 1 1
use contact_7  contact_7_239
timestamp 1624857261
transform 1 0 6041 0 1 3167
box 0 0 1 1
use contact_19  contact_19_239
timestamp 1624857261
transform 1 0 6042 0 1 3172
box 0 0 1 1
use contact_7  contact_7_613
timestamp 1624857261
transform 1 0 6466 0 1 3109
box 0 0 1 1
use contact_19  contact_19_613
timestamp 1624857261
transform 1 0 6467 0 1 3114
box 0 0 1 1
use contact_7  contact_7_611
timestamp 1624857261
transform 1 0 6898 0 1 3109
box 0 0 1 1
use contact_19  contact_19_611
timestamp 1624857261
transform 1 0 6899 0 1 3114
box 0 0 1 1
use contact_7  contact_7_238
timestamp 1624857261
transform 1 0 7280 0 1 3123
box 0 0 1 1
use contact_19  contact_19_238
timestamp 1624857261
transform 1 0 7281 0 1 3128
box 0 0 1 1
use and3_dec  and3_dec_119
timestamp 1624857261
transform 1 0 5803 0 1 3160
box 0 -60 2072 490
use contact_7  contact_7_630
timestamp 1624857261
transform 1 0 7676 0 1 753
box 0 0 1 1
use contact_19  contact_19_630
timestamp 1624857261
transform 1 0 7677 0 1 758
box 0 0 1 1
use contact_7  contact_7_633
timestamp 1624857261
transform 1 0 7676 0 1 358
box 0 0 1 1
use contact_19  contact_19_633
timestamp 1624857261
transform 1 0 7677 0 1 363
box 0 0 1 1
use contact_7  contact_7_624
timestamp 1624857261
transform 1 0 7676 0 1 1543
box 0 0 1 1
use contact_19  contact_19_624
timestamp 1624857261
transform 1 0 7677 0 1 1548
box 0 0 1 1
use contact_7  contact_7_627
timestamp 1624857261
transform 1 0 7676 0 1 1148
box 0 0 1 1
use contact_19  contact_19_627
timestamp 1624857261
transform 1 0 7677 0 1 1153
box 0 0 1 1
use contact_7  contact_7_618
timestamp 1624857261
transform 1 0 7676 0 1 2333
box 0 0 1 1
use contact_19  contact_19_618
timestamp 1624857261
transform 1 0 7677 0 1 2338
box 0 0 1 1
use contact_7  contact_7_621
timestamp 1624857261
transform 1 0 7676 0 1 1938
box 0 0 1 1
use contact_19  contact_19_621
timestamp 1624857261
transform 1 0 7677 0 1 1943
box 0 0 1 1
use contact_7  contact_7_612
timestamp 1624857261
transform 1 0 7676 0 1 3123
box 0 0 1 1
use contact_19  contact_19_612
timestamp 1624857261
transform 1 0 7677 0 1 3128
box 0 0 1 1
use contact_7  contact_7_615
timestamp 1624857261
transform 1 0 7676 0 1 2728
box 0 0 1 1
use contact_19  contact_19_615
timestamp 1624857261
transform 1 0 7677 0 1 2733
box 0 0 1 1
use hierarchical_predecode3x8  hierarchical_predecode3x8_0
timestamp 1624857261
transform 1 0 607 0 1 4740
box 61 -60 3854 3220
use contact_14  contact_14_18
timestamp 1624857261
transform 1 0 672 0 1 4877
box 0 0 1 1
use contact_17  contact_17_386
timestamp 1624857261
transform 1 0 320 0 1 4881
box 0 0 1 1
use contact_14  contact_14_17
timestamp 1624857261
transform 1 0 752 0 1 5327
box 0 0 1 1
use contact_17  contact_17_385
timestamp 1624857261
transform 1 0 400 0 1 5331
box 0 0 1 1
use contact_14  contact_14_16
timestamp 1624857261
transform 1 0 832 0 1 5667
box 0 0 1 1
use contact_17  contact_17_384
timestamp 1624857261
transform 1 0 480 0 1 5671
box 0 0 1 1
use contact_14  contact_14_9
timestamp 1624857261
transform 1 0 4414 0 1 3247
box 0 0 1 1
use contact_19  contact_19_644
timestamp 1624857261
transform 1 0 4411 0 1 3248
box 0 0 1 1
use contact_17  contact_17_358
timestamp 1624857261
transform 1 0 4984 0 1 3324
box 0 0 1 1
use contact_17  contact_17_357
timestamp 1624857261
transform 1 0 5144 0 1 3414
box 0 0 1 1
use contact_17  contact_17_354
timestamp 1624857261
transform 1 0 5144 0 1 3638
box 0 0 1 1
use contact_17  contact_17_355
timestamp 1624857261
transform 1 0 4984 0 1 3728
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1624857261
transform 1 0 5065 0 1 3523
box 0 0 1 1
use contact_7  contact_7_237
timestamp 1624857261
transform 1 0 6041 0 1 3541
box 0 0 1 1
use contact_19  contact_19_237
timestamp 1624857261
transform 1 0 6042 0 1 3546
box 0 0 1 1
use contact_7  contact_7_610
timestamp 1624857261
transform 1 0 6466 0 1 3541
box 0 0 1 1
use contact_19  contact_19_610
timestamp 1624857261
transform 1 0 6467 0 1 3546
box 0 0 1 1
use contact_7  contact_7_608
timestamp 1624857261
transform 1 0 6898 0 1 3541
box 0 0 1 1
use contact_19  contact_19_608
timestamp 1624857261
transform 1 0 6899 0 1 3546
box 0 0 1 1
use contact_7  contact_7_236
timestamp 1624857261
transform 1 0 7280 0 1 3518
box 0 0 1 1
use contact_19  contact_19_236
timestamp 1624857261
transform 1 0 7281 0 1 3523
box 0 0 1 1
use and3_dec  and3_dec_118
timestamp 1624857261
transform 1 0 5803 0 -1 3950
box 0 -60 2072 490
use contact_19  contact_19_643
timestamp 1624857261
transform 1 0 4411 0 1 3798
box 0 0 1 1
use contact_14  contact_14_8
timestamp 1624857261
transform 1 0 4414 0 1 3797
box 0 0 1 1
use contact_17  contact_17_353
timestamp 1624857261
transform 1 0 4664 0 1 4002
box 0 0 1 1
use contact_17  contact_17_356
timestamp 1624857261
transform 1 0 4584 0 1 3840
box 0 0 1 1
use contact_7  contact_7_235
timestamp 1624857261
transform 1 0 6041 0 1 3957
box 0 0 1 1
use contact_19  contact_19_235
timestamp 1624857261
transform 1 0 6042 0 1 3962
box 0 0 1 1
use contact_7  contact_7_607
timestamp 1624857261
transform 1 0 6466 0 1 3899
box 0 0 1 1
use contact_19  contact_19_607
timestamp 1624857261
transform 1 0 6467 0 1 3904
box 0 0 1 1
use contact_7  contact_7_605
timestamp 1624857261
transform 1 0 6898 0 1 3899
box 0 0 1 1
use contact_19  contact_19_605
timestamp 1624857261
transform 1 0 6899 0 1 3904
box 0 0 1 1
use contact_7  contact_7_234
timestamp 1624857261
transform 1 0 7280 0 1 3913
box 0 0 1 1
use contact_19  contact_19_234
timestamp 1624857261
transform 1 0 7281 0 1 3918
box 0 0 1 1
use contact_17  contact_17_352
timestamp 1624857261
transform 1 0 4984 0 1 4114
box 0 0 1 1
use contact_17  contact_17_351
timestamp 1624857261
transform 1 0 5144 0 1 4204
box 0 0 1 1
use contact_19  contact_19_232
timestamp 1624857261
transform 1 0 7281 0 1 4313
box 0 0 1 1
use contact_7  contact_7_232
timestamp 1624857261
transform 1 0 7280 0 1 4308
box 0 0 1 1
use and3_dec  and3_dec_117
timestamp 1624857261
transform 1 0 5803 0 1 3950
box 0 -60 2072 490
use and3_dec  and3_dec_116
timestamp 1624857261
transform 1 0 5803 0 -1 4740
box 0 -60 2072 490
use contact_17  contact_17_349
timestamp 1624857261
transform 1 0 4984 0 1 4518
box 0 0 1 1
use contact_17  contact_17_348
timestamp 1624857261
transform 1 0 5144 0 1 4428
box 0 0 1 1
use contact_19  contact_19_604
timestamp 1624857261
transform 1 0 6467 0 1 4336
box 0 0 1 1
use contact_7  contact_7_604
timestamp 1624857261
transform 1 0 6466 0 1 4331
box 0 0 1 1
use contact_19  contact_19_602
timestamp 1624857261
transform 1 0 6899 0 1 4336
box 0 0 1 1
use contact_7  contact_7_602
timestamp 1624857261
transform 1 0 6898 0 1 4331
box 0 0 1 1
use contact_19  contact_19_233
timestamp 1624857261
transform 1 0 6042 0 1 4336
box 0 0 1 1
use contact_7  contact_7_233
timestamp 1624857261
transform 1 0 6041 0 1 4331
box 0 0 1 1
use contact_17  contact_17_347
timestamp 1624857261
transform 1 0 4504 0 1 4792
box 0 0 1 1
use contact_19  contact_19_642
timestamp 1624857261
transform 1 0 4411 0 1 4828
box 0 0 1 1
use contact_14  contact_14_7
timestamp 1624857261
transform 1 0 4414 0 1 4827
box 0 0 1 1
use contact_17  contact_17_350
timestamp 1624857261
transform 1 0 4744 0 1 4630
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1624857261
transform 1 0 5145 0 1 4708
box 0 0 1 1
use contact_7  contact_7_231
timestamp 1624857261
transform 1 0 6041 0 1 4747
box 0 0 1 1
use contact_19  contact_19_231
timestamp 1624857261
transform 1 0 6042 0 1 4752
box 0 0 1 1
use contact_7  contact_7_601
timestamp 1624857261
transform 1 0 6466 0 1 4689
box 0 0 1 1
use contact_19  contact_19_601
timestamp 1624857261
transform 1 0 6467 0 1 4694
box 0 0 1 1
use contact_7  contact_7_599
timestamp 1624857261
transform 1 0 6898 0 1 4689
box 0 0 1 1
use contact_19  contact_19_599
timestamp 1624857261
transform 1 0 6899 0 1 4694
box 0 0 1 1
use contact_7  contact_7_230
timestamp 1624857261
transform 1 0 7280 0 1 4703
box 0 0 1 1
use contact_19  contact_19_230
timestamp 1624857261
transform 1 0 7281 0 1 4708
box 0 0 1 1
use and3_dec  and3_dec_115
timestamp 1624857261
transform 1 0 5803 0 1 4740
box 0 -60 2072 490
use contact_17  contact_17_345
timestamp 1624857261
transform 1 0 5144 0 1 4994
box 0 0 1 1
use contact_17  contact_17_346
timestamp 1624857261
transform 1 0 5064 0 1 4904
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1624857261
transform 1 0 5225 0 1 5103
box 0 0 1 1
use contact_7  contact_7_229
timestamp 1624857261
transform 1 0 6041 0 1 5121
box 0 0 1 1
use contact_19  contact_19_229
timestamp 1624857261
transform 1 0 6042 0 1 5126
box 0 0 1 1
use contact_7  contact_7_598
timestamp 1624857261
transform 1 0 6466 0 1 5121
box 0 0 1 1
use contact_19  contact_19_598
timestamp 1624857261
transform 1 0 6467 0 1 5126
box 0 0 1 1
use contact_7  contact_7_596
timestamp 1624857261
transform 1 0 6898 0 1 5121
box 0 0 1 1
use contact_19  contact_19_596
timestamp 1624857261
transform 1 0 6899 0 1 5126
box 0 0 1 1
use contact_7  contact_7_228
timestamp 1624857261
transform 1 0 7280 0 1 5098
box 0 0 1 1
use contact_19  contact_19_228
timestamp 1624857261
transform 1 0 7281 0 1 5103
box 0 0 1 1
use contact_14  contact_14_6
timestamp 1624857261
transform 1 0 4414 0 1 5377
box 0 0 1 1
use contact_19  contact_19_641
timestamp 1624857261
transform 1 0 4411 0 1 5378
box 0 0 1 1
use contact_17  contact_17_344
timestamp 1624857261
transform 1 0 4584 0 1 5420
box 0 0 1 1
use contact_17  contact_17_343
timestamp 1624857261
transform 1 0 5064 0 1 5308
box 0 0 1 1
use contact_17  contact_17_342
timestamp 1624857261
transform 1 0 5144 0 1 5218
box 0 0 1 1
use and3_dec  and3_dec_114
timestamp 1624857261
transform 1 0 5803 0 -1 5530
box 0 -60 2072 490
use contact_17  contact_17_341
timestamp 1624857261
transform 1 0 4664 0 1 5582
box 0 0 1 1
use contact_19  contact_19_640
timestamp 1624857261
transform 1 0 4411 0 1 5618
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1624857261
transform 1 0 4414 0 1 5617
box 0 0 1 1
use contact_17  contact_17_340
timestamp 1624857261
transform 1 0 5064 0 1 5694
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1624857261
transform 1 0 5305 0 1 5498
box 0 0 1 1
use contact_7  contact_7_227
timestamp 1624857261
transform 1 0 6041 0 1 5537
box 0 0 1 1
use contact_19  contact_19_227
timestamp 1624857261
transform 1 0 6042 0 1 5542
box 0 0 1 1
use contact_7  contact_7_595
timestamp 1624857261
transform 1 0 6466 0 1 5479
box 0 0 1 1
use contact_19  contact_19_595
timestamp 1624857261
transform 1 0 6467 0 1 5484
box 0 0 1 1
use contact_7  contact_7_593
timestamp 1624857261
transform 1 0 6898 0 1 5479
box 0 0 1 1
use contact_19  contact_19_593
timestamp 1624857261
transform 1 0 6899 0 1 5484
box 0 0 1 1
use contact_7  contact_7_226
timestamp 1624857261
transform 1 0 7280 0 1 5493
box 0 0 1 1
use contact_19  contact_19_226
timestamp 1624857261
transform 1 0 7281 0 1 5498
box 0 0 1 1
use contact_17  contact_17_339
timestamp 1624857261
transform 1 0 5144 0 1 5784
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1624857261
transform 1 0 5385 0 1 5893
box 0 0 1 1
use contact_7  contact_7_225
timestamp 1624857261
transform 1 0 6041 0 1 5911
box 0 0 1 1
use contact_19  contact_19_225
timestamp 1624857261
transform 1 0 6042 0 1 5916
box 0 0 1 1
use contact_7  contact_7_592
timestamp 1624857261
transform 1 0 6466 0 1 5911
box 0 0 1 1
use contact_19  contact_19_592
timestamp 1624857261
transform 1 0 6467 0 1 5916
box 0 0 1 1
use contact_7  contact_7_590
timestamp 1624857261
transform 1 0 6898 0 1 5911
box 0 0 1 1
use contact_19  contact_19_590
timestamp 1624857261
transform 1 0 6899 0 1 5916
box 0 0 1 1
use contact_7  contact_7_224
timestamp 1624857261
transform 1 0 7280 0 1 5888
box 0 0 1 1
use contact_19  contact_19_224
timestamp 1624857261
transform 1 0 7281 0 1 5893
box 0 0 1 1
use and3_dec  and3_dec_113
timestamp 1624857261
transform 1 0 5803 0 1 5530
box 0 -60 2072 490
use and3_dec  and3_dec_112
timestamp 1624857261
transform 1 0 5803 0 -1 6320
box 0 -60 2072 490
use contact_14  contact_14_4
timestamp 1624857261
transform 1 0 4414 0 1 6167
box 0 0 1 1
use contact_19  contact_19_639
timestamp 1624857261
transform 1 0 4411 0 1 6168
box 0 0 1 1
use contact_17  contact_17_338
timestamp 1624857261
transform 1 0 4744 0 1 6210
box 0 0 1 1
use contact_17  contact_17_337
timestamp 1624857261
transform 1 0 5064 0 1 6098
box 0 0 1 1
use contact_17  contact_17_336
timestamp 1624857261
transform 1 0 5144 0 1 6008
box 0 0 1 1
use contact_17  contact_17_335
timestamp 1624857261
transform 1 0 4504 0 1 6372
box 0 0 1 1
use contact_19  contact_19_638
timestamp 1624857261
transform 1 0 4411 0 1 6408
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1624857261
transform 1 0 4414 0 1 6407
box 0 0 1 1
use contact_17  contact_17_334
timestamp 1624857261
transform 1 0 4824 0 1 6484
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1624857261
transform 1 0 5465 0 1 6288
box 0 0 1 1
use contact_7  contact_7_223
timestamp 1624857261
transform 1 0 6041 0 1 6327
box 0 0 1 1
use contact_19  contact_19_223
timestamp 1624857261
transform 1 0 6042 0 1 6332
box 0 0 1 1
use contact_7  contact_7_589
timestamp 1624857261
transform 1 0 6466 0 1 6269
box 0 0 1 1
use contact_19  contact_19_589
timestamp 1624857261
transform 1 0 6467 0 1 6274
box 0 0 1 1
use contact_7  contact_7_587
timestamp 1624857261
transform 1 0 6898 0 1 6269
box 0 0 1 1
use contact_19  contact_19_587
timestamp 1624857261
transform 1 0 6899 0 1 6274
box 0 0 1 1
use contact_7  contact_7_222
timestamp 1624857261
transform 1 0 7280 0 1 6283
box 0 0 1 1
use contact_19  contact_19_222
timestamp 1624857261
transform 1 0 7281 0 1 6288
box 0 0 1 1
use and3_dec  and3_dec_111
timestamp 1624857261
transform 1 0 5803 0 1 6320
box 0 -60 2072 490
use contact_7  contact_7_606
timestamp 1624857261
transform 1 0 7676 0 1 3913
box 0 0 1 1
use contact_19  contact_19_606
timestamp 1624857261
transform 1 0 7677 0 1 3918
box 0 0 1 1
use contact_7  contact_7_609
timestamp 1624857261
transform 1 0 7676 0 1 3518
box 0 0 1 1
use contact_19  contact_19_609
timestamp 1624857261
transform 1 0 7677 0 1 3523
box 0 0 1 1
use contact_7  contact_7_600
timestamp 1624857261
transform 1 0 7676 0 1 4703
box 0 0 1 1
use contact_19  contact_19_600
timestamp 1624857261
transform 1 0 7677 0 1 4708
box 0 0 1 1
use contact_7  contact_7_603
timestamp 1624857261
transform 1 0 7676 0 1 4308
box 0 0 1 1
use contact_19  contact_19_603
timestamp 1624857261
transform 1 0 7677 0 1 4313
box 0 0 1 1
use contact_7  contact_7_594
timestamp 1624857261
transform 1 0 7676 0 1 5493
box 0 0 1 1
use contact_19  contact_19_594
timestamp 1624857261
transform 1 0 7677 0 1 5498
box 0 0 1 1
use contact_7  contact_7_597
timestamp 1624857261
transform 1 0 7676 0 1 5098
box 0 0 1 1
use contact_19  contact_19_597
timestamp 1624857261
transform 1 0 7677 0 1 5103
box 0 0 1 1
use contact_7  contact_7_588
timestamp 1624857261
transform 1 0 7676 0 1 6283
box 0 0 1 1
use contact_19  contact_19_588
timestamp 1624857261
transform 1 0 7677 0 1 6288
box 0 0 1 1
use contact_7  contact_7_591
timestamp 1624857261
transform 1 0 7676 0 1 5888
box 0 0 1 1
use contact_19  contact_19_591
timestamp 1624857261
transform 1 0 7677 0 1 5893
box 0 0 1 1
use contact_17  contact_17_333
timestamp 1624857261
transform 1 0 5224 0 1 6574
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1624857261
transform 1 0 5545 0 1 6683
box 0 0 1 1
use contact_7  contact_7_221
timestamp 1624857261
transform 1 0 6041 0 1 6701
box 0 0 1 1
use contact_19  contact_19_221
timestamp 1624857261
transform 1 0 6042 0 1 6706
box 0 0 1 1
use contact_7  contact_7_586
timestamp 1624857261
transform 1 0 6466 0 1 6701
box 0 0 1 1
use contact_19  contact_19_586
timestamp 1624857261
transform 1 0 6467 0 1 6706
box 0 0 1 1
use contact_7  contact_7_584
timestamp 1624857261
transform 1 0 6898 0 1 6701
box 0 0 1 1
use contact_19  contact_19_584
timestamp 1624857261
transform 1 0 6899 0 1 6706
box 0 0 1 1
use contact_7  contact_7_220
timestamp 1624857261
transform 1 0 7280 0 1 6678
box 0 0 1 1
use contact_19  contact_19_220
timestamp 1624857261
transform 1 0 7281 0 1 6683
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1624857261
transform 1 0 4414 0 1 6957
box 0 0 1 1
use contact_19  contact_19_637
timestamp 1624857261
transform 1 0 4411 0 1 6958
box 0 0 1 1
use contact_17  contact_17_332
timestamp 1624857261
transform 1 0 4584 0 1 7000
box 0 0 1 1
use contact_17  contact_17_331
timestamp 1624857261
transform 1 0 4824 0 1 6888
box 0 0 1 1
use contact_17  contact_17_330
timestamp 1624857261
transform 1 0 5224 0 1 6798
box 0 0 1 1
use and3_dec  and3_dec_110
timestamp 1624857261
transform 1 0 5803 0 -1 7110
box 0 -60 2072 490
use and3_dec  and3_dec_109
timestamp 1624857261
transform 1 0 5803 0 1 7110
box 0 -60 2072 490
use contact_17  contact_17_329
timestamp 1624857261
transform 1 0 4664 0 1 7162
box 0 0 1 1
use contact_19  contact_19_636
timestamp 1624857261
transform 1 0 4411 0 1 7198
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1624857261
transform 1 0 4414 0 1 7197
box 0 0 1 1
use contact_17  contact_17_328
timestamp 1624857261
transform 1 0 4824 0 1 7274
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1624857261
transform 1 0 5625 0 1 7078
box 0 0 1 1
use contact_7  contact_7_219
timestamp 1624857261
transform 1 0 6041 0 1 7117
box 0 0 1 1
use contact_19  contact_19_219
timestamp 1624857261
transform 1 0 6042 0 1 7122
box 0 0 1 1
use contact_7  contact_7_583
timestamp 1624857261
transform 1 0 6466 0 1 7059
box 0 0 1 1
use contact_19  contact_19_583
timestamp 1624857261
transform 1 0 6467 0 1 7064
box 0 0 1 1
use contact_7  contact_7_581
timestamp 1624857261
transform 1 0 6898 0 1 7059
box 0 0 1 1
use contact_19  contact_19_581
timestamp 1624857261
transform 1 0 6899 0 1 7064
box 0 0 1 1
use contact_7  contact_7_218
timestamp 1624857261
transform 1 0 7280 0 1 7073
box 0 0 1 1
use contact_19  contact_19_218
timestamp 1624857261
transform 1 0 7281 0 1 7078
box 0 0 1 1
use contact_17  contact_17_324
timestamp 1624857261
transform 1 0 5224 0 1 7588
box 0 0 1 1
use contact_17  contact_17_327
timestamp 1624857261
transform 1 0 5224 0 1 7364
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1624857261
transform 1 0 5705 0 1 7473
box 0 0 1 1
use contact_7  contact_7_217
timestamp 1624857261
transform 1 0 6041 0 1 7491
box 0 0 1 1
use contact_19  contact_19_217
timestamp 1624857261
transform 1 0 6042 0 1 7496
box 0 0 1 1
use contact_7  contact_7_580
timestamp 1624857261
transform 1 0 6466 0 1 7491
box 0 0 1 1
use contact_19  contact_19_580
timestamp 1624857261
transform 1 0 6467 0 1 7496
box 0 0 1 1
use contact_7  contact_7_578
timestamp 1624857261
transform 1 0 6898 0 1 7491
box 0 0 1 1
use contact_19  contact_19_578
timestamp 1624857261
transform 1 0 6899 0 1 7496
box 0 0 1 1
use contact_7  contact_7_216
timestamp 1624857261
transform 1 0 7280 0 1 7468
box 0 0 1 1
use contact_19  contact_19_216
timestamp 1624857261
transform 1 0 7281 0 1 7473
box 0 0 1 1
use and3_dec  and3_dec_108
timestamp 1624857261
transform 1 0 5803 0 -1 7900
box 0 -60 2072 490
use contact_19  contact_19_635
timestamp 1624857261
transform 1 0 4411 0 1 7748
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1624857261
transform 1 0 4414 0 1 7747
box 0 0 1 1
use contact_17  contact_17_325
timestamp 1624857261
transform 1 0 4824 0 1 7678
box 0 0 1 1
use contact_17  contact_17_326
timestamp 1624857261
transform 1 0 4744 0 1 7790
box 0 0 1 1
use contact_7  contact_7_577
timestamp 1624857261
transform 1 0 6466 0 1 7849
box 0 0 1 1
use contact_19  contact_19_577
timestamp 1624857261
transform 1 0 6467 0 1 7854
box 0 0 1 1
use contact_7  contact_7_575
timestamp 1624857261
transform 1 0 6898 0 1 7849
box 0 0 1 1
use contact_19  contact_19_575
timestamp 1624857261
transform 1 0 6899 0 1 7854
box 0 0 1 1
use contact_7  contact_7_214
timestamp 1624857261
transform 1 0 7280 0 1 7863
box 0 0 1 1
use contact_19  contact_19_214
timestamp 1624857261
transform 1 0 7281 0 1 7868
box 0 0 1 1
use contact_17  contact_17_323
timestamp 1624857261
transform 1 0 4504 0 1 7952
box 0 0 1 1
use contact_17  contact_17_322
timestamp 1624857261
transform 1 0 4904 0 1 8064
box 0 0 1 1
use contact_17  contact_17_321
timestamp 1624857261
transform 1 0 5224 0 1 8154
box 0 0 1 1
use contact_19  contact_19_215
timestamp 1624857261
transform 1 0 6042 0 1 7912
box 0 0 1 1
use contact_7  contact_7_215
timestamp 1624857261
transform 1 0 6041 0 1 7907
box 0 0 1 1
use and3_dec  and3_dec_107
timestamp 1624857261
transform 1 0 5803 0 1 7900
box 0 -60 2072 490
use contact_17  contact_17_318
timestamp 1624857261
transform 1 0 5224 0 1 8378
box 0 0 1 1
use contact_19  contact_19_574
timestamp 1624857261
transform 1 0 6467 0 1 8286
box 0 0 1 1
use contact_7  contact_7_574
timestamp 1624857261
transform 1 0 6466 0 1 8281
box 0 0 1 1
use contact_19  contact_19_572
timestamp 1624857261
transform 1 0 6899 0 1 8286
box 0 0 1 1
use contact_7  contact_7_572
timestamp 1624857261
transform 1 0 6898 0 1 8281
box 0 0 1 1
use contact_19  contact_19_213
timestamp 1624857261
transform 1 0 6042 0 1 8286
box 0 0 1 1
use contact_7  contact_7_213
timestamp 1624857261
transform 1 0 6041 0 1 8281
box 0 0 1 1
use contact_19  contact_19_212
timestamp 1624857261
transform 1 0 7281 0 1 8263
box 0 0 1 1
use contact_7  contact_7_212
timestamp 1624857261
transform 1 0 7280 0 1 8258
box 0 0 1 1
use contact_17  contact_17_319
timestamp 1624857261
transform 1 0 4904 0 1 8468
box 0 0 1 1
use contact_17  contact_17_320
timestamp 1624857261
transform 1 0 4584 0 1 8580
box 0 0 1 1
use contact_7  contact_7_211
timestamp 1624857261
transform 1 0 6041 0 1 8697
box 0 0 1 1
use contact_19  contact_19_211
timestamp 1624857261
transform 1 0 6042 0 1 8702
box 0 0 1 1
use contact_7  contact_7_571
timestamp 1624857261
transform 1 0 6466 0 1 8639
box 0 0 1 1
use contact_19  contact_19_571
timestamp 1624857261
transform 1 0 6467 0 1 8644
box 0 0 1 1
use contact_7  contact_7_569
timestamp 1624857261
transform 1 0 6898 0 1 8639
box 0 0 1 1
use contact_19  contact_19_569
timestamp 1624857261
transform 1 0 6899 0 1 8644
box 0 0 1 1
use contact_7  contact_7_210
timestamp 1624857261
transform 1 0 7280 0 1 8653
box 0 0 1 1
use contact_19  contact_19_210
timestamp 1624857261
transform 1 0 7281 0 1 8658
box 0 0 1 1
use and3_dec  and3_dec_106
timestamp 1624857261
transform 1 0 5803 0 -1 8690
box 0 -60 2072 490
use and3_dec  and3_dec_105
timestamp 1624857261
transform 1 0 5803 0 1 8690
box 0 -60 2072 490
use contact_17  contact_17_317
timestamp 1624857261
transform 1 0 4664 0 1 8742
box 0 0 1 1
use contact_17  contact_17_316
timestamp 1624857261
transform 1 0 4904 0 1 8854
box 0 0 1 1
use contact_17  contact_17_315
timestamp 1624857261
transform 1 0 5224 0 1 8944
box 0 0 1 1
use contact_17  contact_17_312
timestamp 1624857261
transform 1 0 5224 0 1 9168
box 0 0 1 1
use contact_19  contact_19_568
timestamp 1624857261
transform 1 0 6467 0 1 9076
box 0 0 1 1
use contact_7  contact_7_568
timestamp 1624857261
transform 1 0 6466 0 1 9071
box 0 0 1 1
use contact_19  contact_19_566
timestamp 1624857261
transform 1 0 6899 0 1 9076
box 0 0 1 1
use contact_7  contact_7_566
timestamp 1624857261
transform 1 0 6898 0 1 9071
box 0 0 1 1
use contact_19  contact_19_209
timestamp 1624857261
transform 1 0 6042 0 1 9076
box 0 0 1 1
use contact_7  contact_7_209
timestamp 1624857261
transform 1 0 6041 0 1 9071
box 0 0 1 1
use contact_19  contact_19_208
timestamp 1624857261
transform 1 0 7281 0 1 9053
box 0 0 1 1
use contact_7  contact_7_208
timestamp 1624857261
transform 1 0 7280 0 1 9048
box 0 0 1 1
use and3_dec  and3_dec_104
timestamp 1624857261
transform 1 0 5803 0 -1 9480
box 0 -60 2072 490
use contact_17  contact_17_311
timestamp 1624857261
transform 1 0 4504 0 1 9532
box 0 0 1 1
use contact_17  contact_17_314
timestamp 1624857261
transform 1 0 4744 0 1 9370
box 0 0 1 1
use contact_17  contact_17_313
timestamp 1624857261
transform 1 0 4904 0 1 9258
box 0 0 1 1
use contact_7  contact_7_207
timestamp 1624857261
transform 1 0 6041 0 1 9487
box 0 0 1 1
use contact_19  contact_19_207
timestamp 1624857261
transform 1 0 6042 0 1 9492
box 0 0 1 1
use contact_7  contact_7_565
timestamp 1624857261
transform 1 0 6466 0 1 9429
box 0 0 1 1
use contact_19  contact_19_565
timestamp 1624857261
transform 1 0 6467 0 1 9434
box 0 0 1 1
use contact_7  contact_7_563
timestamp 1624857261
transform 1 0 6898 0 1 9429
box 0 0 1 1
use contact_19  contact_19_563
timestamp 1624857261
transform 1 0 6899 0 1 9434
box 0 0 1 1
use contact_7  contact_7_206
timestamp 1624857261
transform 1 0 7280 0 1 9443
box 0 0 1 1
use contact_19  contact_19_206
timestamp 1624857261
transform 1 0 7281 0 1 9448
box 0 0 1 1
use contact_17  contact_17_310
timestamp 1624857261
transform 1 0 4984 0 1 9644
box 0 0 1 1
use contact_17  contact_17_309
timestamp 1624857261
transform 1 0 5224 0 1 9734
box 0 0 1 1
use and3_dec  and3_dec_103
timestamp 1624857261
transform 1 0 5803 0 1 9480
box 0 -60 2072 490
use and3_dec  and3_dec_102
timestamp 1624857261
transform 1 0 5803 0 -1 10270
box 0 -60 2072 490
use contact_7  contact_7_582
timestamp 1624857261
transform 1 0 7676 0 1 7073
box 0 0 1 1
use contact_19  contact_19_582
timestamp 1624857261
transform 1 0 7677 0 1 7078
box 0 0 1 1
use contact_7  contact_7_585
timestamp 1624857261
transform 1 0 7676 0 1 6678
box 0 0 1 1
use contact_19  contact_19_585
timestamp 1624857261
transform 1 0 7677 0 1 6683
box 0 0 1 1
use contact_7  contact_7_573
timestamp 1624857261
transform 1 0 7676 0 1 8258
box 0 0 1 1
use contact_19  contact_19_573
timestamp 1624857261
transform 1 0 7677 0 1 8263
box 0 0 1 1
use contact_7  contact_7_576
timestamp 1624857261
transform 1 0 7676 0 1 7863
box 0 0 1 1
use contact_19  contact_19_576
timestamp 1624857261
transform 1 0 7677 0 1 7868
box 0 0 1 1
use contact_7  contact_7_579
timestamp 1624857261
transform 1 0 7676 0 1 7468
box 0 0 1 1
use contact_19  contact_19_579
timestamp 1624857261
transform 1 0 7677 0 1 7473
box 0 0 1 1
use contact_7  contact_7_567
timestamp 1624857261
transform 1 0 7676 0 1 9048
box 0 0 1 1
use contact_19  contact_19_567
timestamp 1624857261
transform 1 0 7677 0 1 9053
box 0 0 1 1
use contact_7  contact_7_570
timestamp 1624857261
transform 1 0 7676 0 1 8653
box 0 0 1 1
use contact_19  contact_19_570
timestamp 1624857261
transform 1 0 7677 0 1 8658
box 0 0 1 1
use contact_7  contact_7_564
timestamp 1624857261
transform 1 0 7676 0 1 9443
box 0 0 1 1
use contact_19  contact_19_564
timestamp 1624857261
transform 1 0 7677 0 1 9448
box 0 0 1 1
use contact_17  contact_17_306
timestamp 1624857261
transform 1 0 5224 0 1 9958
box 0 0 1 1
use contact_17  contact_17_307
timestamp 1624857261
transform 1 0 4984 0 1 10048
box 0 0 1 1
use contact_7  contact_7_205
timestamp 1624857261
transform 1 0 6041 0 1 9861
box 0 0 1 1
use contact_19  contact_19_205
timestamp 1624857261
transform 1 0 6042 0 1 9866
box 0 0 1 1
use contact_7  contact_7_562
timestamp 1624857261
transform 1 0 6466 0 1 9861
box 0 0 1 1
use contact_19  contact_19_562
timestamp 1624857261
transform 1 0 6467 0 1 9866
box 0 0 1 1
use contact_7  contact_7_560
timestamp 1624857261
transform 1 0 6898 0 1 9861
box 0 0 1 1
use contact_19  contact_19_560
timestamp 1624857261
transform 1 0 6899 0 1 9866
box 0 0 1 1
use contact_7  contact_7_204
timestamp 1624857261
transform 1 0 7280 0 1 9838
box 0 0 1 1
use contact_19  contact_19_204
timestamp 1624857261
transform 1 0 7281 0 1 9843
box 0 0 1 1
use contact_17  contact_17_305
timestamp 1624857261
transform 1 0 4664 0 1 10322
box 0 0 1 1
use contact_17  contact_17_308
timestamp 1624857261
transform 1 0 4584 0 1 10160
box 0 0 1 1
use contact_7  contact_7_203
timestamp 1624857261
transform 1 0 6041 0 1 10277
box 0 0 1 1
use contact_19  contact_19_203
timestamp 1624857261
transform 1 0 6042 0 1 10282
box 0 0 1 1
use contact_7  contact_7_559
timestamp 1624857261
transform 1 0 6466 0 1 10219
box 0 0 1 1
use contact_19  contact_19_559
timestamp 1624857261
transform 1 0 6467 0 1 10224
box 0 0 1 1
use contact_7  contact_7_557
timestamp 1624857261
transform 1 0 6898 0 1 10219
box 0 0 1 1
use contact_19  contact_19_557
timestamp 1624857261
transform 1 0 6899 0 1 10224
box 0 0 1 1
use contact_7  contact_7_202
timestamp 1624857261
transform 1 0 7280 0 1 10233
box 0 0 1 1
use contact_19  contact_19_202
timestamp 1624857261
transform 1 0 7281 0 1 10238
box 0 0 1 1
use and3_dec  and3_dec_101
timestamp 1624857261
transform 1 0 5803 0 1 10270
box 0 -60 2072 490
use contact_17  contact_17_304
timestamp 1624857261
transform 1 0 4984 0 1 10434
box 0 0 1 1
use contact_17  contact_17_303
timestamp 1624857261
transform 1 0 5224 0 1 10524
box 0 0 1 1
use contact_17  contact_17_300
timestamp 1624857261
transform 1 0 5224 0 1 10748
box 0 0 1 1
use contact_17  contact_17_301
timestamp 1624857261
transform 1 0 4984 0 1 10838
box 0 0 1 1
use contact_7  contact_7_201
timestamp 1624857261
transform 1 0 6041 0 1 10651
box 0 0 1 1
use contact_19  contact_19_201
timestamp 1624857261
transform 1 0 6042 0 1 10656
box 0 0 1 1
use contact_7  contact_7_556
timestamp 1624857261
transform 1 0 6466 0 1 10651
box 0 0 1 1
use contact_19  contact_19_556
timestamp 1624857261
transform 1 0 6467 0 1 10656
box 0 0 1 1
use contact_7  contact_7_554
timestamp 1624857261
transform 1 0 6898 0 1 10651
box 0 0 1 1
use contact_19  contact_19_554
timestamp 1624857261
transform 1 0 6899 0 1 10656
box 0 0 1 1
use contact_7  contact_7_200
timestamp 1624857261
transform 1 0 7280 0 1 10628
box 0 0 1 1
use contact_19  contact_19_200
timestamp 1624857261
transform 1 0 7281 0 1 10633
box 0 0 1 1
use and3_dec  and3_dec_100
timestamp 1624857261
transform 1 0 5803 0 -1 11060
box 0 -60 2072 490
use contact_17  contact_17_299
timestamp 1624857261
transform 1 0 4504 0 1 11112
box 0 0 1 1
use contact_17  contact_17_302
timestamp 1624857261
transform 1 0 4744 0 1 10950
box 0 0 1 1
use contact_7  contact_7_199
timestamp 1624857261
transform 1 0 6041 0 1 11067
box 0 0 1 1
use contact_19  contact_19_199
timestamp 1624857261
transform 1 0 6042 0 1 11072
box 0 0 1 1
use contact_7  contact_7_553
timestamp 1624857261
transform 1 0 6466 0 1 11009
box 0 0 1 1
use contact_19  contact_19_553
timestamp 1624857261
transform 1 0 6467 0 1 11014
box 0 0 1 1
use contact_7  contact_7_551
timestamp 1624857261
transform 1 0 6898 0 1 11009
box 0 0 1 1
use contact_19  contact_19_551
timestamp 1624857261
transform 1 0 6899 0 1 11014
box 0 0 1 1
use contact_7  contact_7_198
timestamp 1624857261
transform 1 0 7280 0 1 11023
box 0 0 1 1
use contact_19  contact_19_198
timestamp 1624857261
transform 1 0 7281 0 1 11028
box 0 0 1 1
use contact_17  contact_17_298
timestamp 1624857261
transform 1 0 5064 0 1 11224
box 0 0 1 1
use contact_17  contact_17_297
timestamp 1624857261
transform 1 0 5224 0 1 11314
box 0 0 1 1
use contact_19  contact_19_196
timestamp 1624857261
transform 1 0 7281 0 1 11423
box 0 0 1 1
use contact_7  contact_7_196
timestamp 1624857261
transform 1 0 7280 0 1 11418
box 0 0 1 1
use and3_dec  and3_dec_99
timestamp 1624857261
transform 1 0 5803 0 1 11060
box 0 -60 2072 490
use and3_dec  and3_dec_98
timestamp 1624857261
transform 1 0 5803 0 -1 11850
box 0 -60 2072 490
use contact_17  contact_17_295
timestamp 1624857261
transform 1 0 5064 0 1 11628
box 0 0 1 1
use contact_17  contact_17_294
timestamp 1624857261
transform 1 0 5224 0 1 11538
box 0 0 1 1
use contact_19  contact_19_550
timestamp 1624857261
transform 1 0 6467 0 1 11446
box 0 0 1 1
use contact_7  contact_7_550
timestamp 1624857261
transform 1 0 6466 0 1 11441
box 0 0 1 1
use contact_19  contact_19_548
timestamp 1624857261
transform 1 0 6899 0 1 11446
box 0 0 1 1
use contact_7  contact_7_548
timestamp 1624857261
transform 1 0 6898 0 1 11441
box 0 0 1 1
use contact_19  contact_19_197
timestamp 1624857261
transform 1 0 6042 0 1 11446
box 0 0 1 1
use contact_7  contact_7_197
timestamp 1624857261
transform 1 0 6041 0 1 11441
box 0 0 1 1
use contact_17  contact_17_293
timestamp 1624857261
transform 1 0 4664 0 1 11902
box 0 0 1 1
use contact_17  contact_17_296
timestamp 1624857261
transform 1 0 4584 0 1 11740
box 0 0 1 1
use contact_7  contact_7_195
timestamp 1624857261
transform 1 0 6041 0 1 11857
box 0 0 1 1
use contact_19  contact_19_195
timestamp 1624857261
transform 1 0 6042 0 1 11862
box 0 0 1 1
use contact_7  contact_7_547
timestamp 1624857261
transform 1 0 6466 0 1 11799
box 0 0 1 1
use contact_19  contact_19_547
timestamp 1624857261
transform 1 0 6467 0 1 11804
box 0 0 1 1
use contact_7  contact_7_545
timestamp 1624857261
transform 1 0 6898 0 1 11799
box 0 0 1 1
use contact_19  contact_19_545
timestamp 1624857261
transform 1 0 6899 0 1 11804
box 0 0 1 1
use contact_7  contact_7_194
timestamp 1624857261
transform 1 0 7280 0 1 11813
box 0 0 1 1
use contact_19  contact_19_194
timestamp 1624857261
transform 1 0 7281 0 1 11818
box 0 0 1 1
use and3_dec  and3_dec_97
timestamp 1624857261
transform 1 0 5803 0 1 11850
box 0 -60 2072 490
use contact_17  contact_17_291
timestamp 1624857261
transform 1 0 5224 0 1 12104
box 0 0 1 1
use contact_17  contact_17_292
timestamp 1624857261
transform 1 0 5064 0 1 12014
box 0 0 1 1
use contact_7  contact_7_193
timestamp 1624857261
transform 1 0 6041 0 1 12231
box 0 0 1 1
use contact_19  contact_19_193
timestamp 1624857261
transform 1 0 6042 0 1 12236
box 0 0 1 1
use contact_7  contact_7_544
timestamp 1624857261
transform 1 0 6466 0 1 12231
box 0 0 1 1
use contact_19  contact_19_544
timestamp 1624857261
transform 1 0 6467 0 1 12236
box 0 0 1 1
use contact_7  contact_7_542
timestamp 1624857261
transform 1 0 6898 0 1 12231
box 0 0 1 1
use contact_19  contact_19_542
timestamp 1624857261
transform 1 0 6899 0 1 12236
box 0 0 1 1
use contact_7  contact_7_192
timestamp 1624857261
transform 1 0 7280 0 1 12208
box 0 0 1 1
use contact_19  contact_19_192
timestamp 1624857261
transform 1 0 7281 0 1 12213
box 0 0 1 1
use contact_17  contact_17_290
timestamp 1624857261
transform 1 0 4744 0 1 12530
box 0 0 1 1
use contact_17  contact_17_289
timestamp 1624857261
transform 1 0 5064 0 1 12418
box 0 0 1 1
use contact_17  contact_17_288
timestamp 1624857261
transform 1 0 5224 0 1 12328
box 0 0 1 1
use and3_dec  and3_dec_96
timestamp 1624857261
transform 1 0 5803 0 -1 12640
box 0 -60 2072 490
use contact_17  contact_17_287
timestamp 1624857261
transform 1 0 4504 0 1 12692
box 0 0 1 1
use contact_17  contact_17_286
timestamp 1624857261
transform 1 0 4824 0 1 12804
box 0 0 1 1
use contact_7  contact_7_191
timestamp 1624857261
transform 1 0 6041 0 1 12647
box 0 0 1 1
use contact_19  contact_19_191
timestamp 1624857261
transform 1 0 6042 0 1 12652
box 0 0 1 1
use contact_7  contact_7_541
timestamp 1624857261
transform 1 0 6466 0 1 12589
box 0 0 1 1
use contact_19  contact_19_541
timestamp 1624857261
transform 1 0 6467 0 1 12594
box 0 0 1 1
use contact_7  contact_7_539
timestamp 1624857261
transform 1 0 6898 0 1 12589
box 0 0 1 1
use contact_19  contact_19_539
timestamp 1624857261
transform 1 0 6899 0 1 12594
box 0 0 1 1
use contact_7  contact_7_190
timestamp 1624857261
transform 1 0 7280 0 1 12603
box 0 0 1 1
use contact_19  contact_19_190
timestamp 1624857261
transform 1 0 7281 0 1 12608
box 0 0 1 1
use contact_17  contact_17_285
timestamp 1624857261
transform 1 0 5304 0 1 12894
box 0 0 1 1
use contact_19  contact_19_538
timestamp 1624857261
transform 1 0 6467 0 1 13026
box 0 0 1 1
use contact_7  contact_7_538
timestamp 1624857261
transform 1 0 6466 0 1 13021
box 0 0 1 1
use contact_19  contact_19_536
timestamp 1624857261
transform 1 0 6899 0 1 13026
box 0 0 1 1
use contact_7  contact_7_536
timestamp 1624857261
transform 1 0 6898 0 1 13021
box 0 0 1 1
use contact_19  contact_19_189
timestamp 1624857261
transform 1 0 6042 0 1 13026
box 0 0 1 1
use contact_7  contact_7_189
timestamp 1624857261
transform 1 0 6041 0 1 13021
box 0 0 1 1
use contact_19  contact_19_188
timestamp 1624857261
transform 1 0 7281 0 1 13003
box 0 0 1 1
use contact_7  contact_7_188
timestamp 1624857261
transform 1 0 7280 0 1 12998
box 0 0 1 1
use and3_dec  and3_dec_95
timestamp 1624857261
transform 1 0 5803 0 1 12640
box 0 -60 2072 490
use and3_dec  and3_dec_94
timestamp 1624857261
transform 1 0 5803 0 -1 13430
box 0 -60 2072 490
use contact_7  contact_7_558
timestamp 1624857261
transform 1 0 7676 0 1 10233
box 0 0 1 1
use contact_19  contact_19_558
timestamp 1624857261
transform 1 0 7677 0 1 10238
box 0 0 1 1
use contact_7  contact_7_561
timestamp 1624857261
transform 1 0 7676 0 1 9838
box 0 0 1 1
use contact_19  contact_19_561
timestamp 1624857261
transform 1 0 7677 0 1 9843
box 0 0 1 1
use contact_7  contact_7_549
timestamp 1624857261
transform 1 0 7676 0 1 11418
box 0 0 1 1
use contact_19  contact_19_549
timestamp 1624857261
transform 1 0 7677 0 1 11423
box 0 0 1 1
use contact_7  contact_7_552
timestamp 1624857261
transform 1 0 7676 0 1 11023
box 0 0 1 1
use contact_19  contact_19_552
timestamp 1624857261
transform 1 0 7677 0 1 11028
box 0 0 1 1
use contact_7  contact_7_555
timestamp 1624857261
transform 1 0 7676 0 1 10628
box 0 0 1 1
use contact_19  contact_19_555
timestamp 1624857261
transform 1 0 7677 0 1 10633
box 0 0 1 1
use contact_7  contact_7_543
timestamp 1624857261
transform 1 0 7676 0 1 12208
box 0 0 1 1
use contact_19  contact_19_543
timestamp 1624857261
transform 1 0 7677 0 1 12213
box 0 0 1 1
use contact_7  contact_7_546
timestamp 1624857261
transform 1 0 7676 0 1 11813
box 0 0 1 1
use contact_19  contact_19_546
timestamp 1624857261
transform 1 0 7677 0 1 11818
box 0 0 1 1
use contact_7  contact_7_537
timestamp 1624857261
transform 1 0 7676 0 1 12998
box 0 0 1 1
use contact_19  contact_19_537
timestamp 1624857261
transform 1 0 7677 0 1 13003
box 0 0 1 1
use contact_7  contact_7_540
timestamp 1624857261
transform 1 0 7676 0 1 12603
box 0 0 1 1
use contact_19  contact_19_540
timestamp 1624857261
transform 1 0 7677 0 1 12608
box 0 0 1 1
use contact_17  contact_17_284
timestamp 1624857261
transform 1 0 4584 0 1 13320
box 0 0 1 1
use contact_17  contact_17_283
timestamp 1624857261
transform 1 0 4824 0 1 13208
box 0 0 1 1
use contact_17  contact_17_282
timestamp 1624857261
transform 1 0 5304 0 1 13118
box 0 0 1 1
use contact_17  contact_17_280
timestamp 1624857261
transform 1 0 4824 0 1 13594
box 0 0 1 1
use contact_17  contact_17_281
timestamp 1624857261
transform 1 0 4664 0 1 13482
box 0 0 1 1
use contact_7  contact_7_187
timestamp 1624857261
transform 1 0 6041 0 1 13437
box 0 0 1 1
use contact_19  contact_19_187
timestamp 1624857261
transform 1 0 6042 0 1 13442
box 0 0 1 1
use contact_7  contact_7_535
timestamp 1624857261
transform 1 0 6466 0 1 13379
box 0 0 1 1
use contact_19  contact_19_535
timestamp 1624857261
transform 1 0 6467 0 1 13384
box 0 0 1 1
use contact_7  contact_7_533
timestamp 1624857261
transform 1 0 6898 0 1 13379
box 0 0 1 1
use contact_19  contact_19_533
timestamp 1624857261
transform 1 0 6899 0 1 13384
box 0 0 1 1
use contact_7  contact_7_186
timestamp 1624857261
transform 1 0 7280 0 1 13393
box 0 0 1 1
use contact_19  contact_19_186
timestamp 1624857261
transform 1 0 7281 0 1 13398
box 0 0 1 1
use and3_dec  and3_dec_93
timestamp 1624857261
transform 1 0 5803 0 1 13430
box 0 -60 2072 490
use contact_17  contact_17_279
timestamp 1624857261
transform 1 0 5304 0 1 13684
box 0 0 1 1
use contact_19  contact_19_532
timestamp 1624857261
transform 1 0 6467 0 1 13816
box 0 0 1 1
use contact_7  contact_7_532
timestamp 1624857261
transform 1 0 6466 0 1 13811
box 0 0 1 1
use contact_19  contact_19_530
timestamp 1624857261
transform 1 0 6899 0 1 13816
box 0 0 1 1
use contact_7  contact_7_530
timestamp 1624857261
transform 1 0 6898 0 1 13811
box 0 0 1 1
use contact_19  contact_19_185
timestamp 1624857261
transform 1 0 6042 0 1 13816
box 0 0 1 1
use contact_7  contact_7_185
timestamp 1624857261
transform 1 0 6041 0 1 13811
box 0 0 1 1
use contact_19  contact_19_184
timestamp 1624857261
transform 1 0 7281 0 1 13793
box 0 0 1 1
use contact_7  contact_7_184
timestamp 1624857261
transform 1 0 7280 0 1 13788
box 0 0 1 1
use contact_17  contact_17_278
timestamp 1624857261
transform 1 0 4744 0 1 14110
box 0 0 1 1
use contact_17  contact_17_277
timestamp 1624857261
transform 1 0 4824 0 1 13998
box 0 0 1 1
use contact_17  contact_17_276
timestamp 1624857261
transform 1 0 5304 0 1 13908
box 0 0 1 1
use and3_dec  and3_dec_92
timestamp 1624857261
transform 1 0 5803 0 -1 14220
box 0 -60 2072 490
use and3_dec  and3_dec_91
timestamp 1624857261
transform 1 0 5803 0 1 14220
box 0 -60 2072 490
use contact_17  contact_17_275
timestamp 1624857261
transform 1 0 4504 0 1 14272
box 0 0 1 1
use contact_17  contact_17_274
timestamp 1624857261
transform 1 0 4904 0 1 14384
box 0 0 1 1
use contact_7  contact_7_183
timestamp 1624857261
transform 1 0 6041 0 1 14227
box 0 0 1 1
use contact_19  contact_19_183
timestamp 1624857261
transform 1 0 6042 0 1 14232
box 0 0 1 1
use contact_7  contact_7_529
timestamp 1624857261
transform 1 0 6466 0 1 14169
box 0 0 1 1
use contact_19  contact_19_529
timestamp 1624857261
transform 1 0 6467 0 1 14174
box 0 0 1 1
use contact_7  contact_7_527
timestamp 1624857261
transform 1 0 6898 0 1 14169
box 0 0 1 1
use contact_19  contact_19_527
timestamp 1624857261
transform 1 0 6899 0 1 14174
box 0 0 1 1
use contact_7  contact_7_182
timestamp 1624857261
transform 1 0 7280 0 1 14183
box 0 0 1 1
use contact_19  contact_19_182
timestamp 1624857261
transform 1 0 7281 0 1 14188
box 0 0 1 1
use contact_17  contact_17_270
timestamp 1624857261
transform 1 0 5304 0 1 14698
box 0 0 1 1
use contact_17  contact_17_273
timestamp 1624857261
transform 1 0 5304 0 1 14474
box 0 0 1 1
use contact_7  contact_7_181
timestamp 1624857261
transform 1 0 6041 0 1 14601
box 0 0 1 1
use contact_19  contact_19_181
timestamp 1624857261
transform 1 0 6042 0 1 14606
box 0 0 1 1
use contact_7  contact_7_526
timestamp 1624857261
transform 1 0 6466 0 1 14601
box 0 0 1 1
use contact_19  contact_19_526
timestamp 1624857261
transform 1 0 6467 0 1 14606
box 0 0 1 1
use contact_7  contact_7_524
timestamp 1624857261
transform 1 0 6898 0 1 14601
box 0 0 1 1
use contact_19  contact_19_524
timestamp 1624857261
transform 1 0 6899 0 1 14606
box 0 0 1 1
use contact_7  contact_7_180
timestamp 1624857261
transform 1 0 7280 0 1 14578
box 0 0 1 1
use contact_19  contact_19_180
timestamp 1624857261
transform 1 0 7281 0 1 14583
box 0 0 1 1
use and3_dec  and3_dec_90
timestamp 1624857261
transform 1 0 5803 0 -1 15010
box 0 -60 2072 490
use contact_17  contact_17_272
timestamp 1624857261
transform 1 0 4584 0 1 14900
box 0 0 1 1
use contact_17  contact_17_271
timestamp 1624857261
transform 1 0 4904 0 1 14788
box 0 0 1 1
use contact_19  contact_19_523
timestamp 1624857261
transform 1 0 6467 0 1 14964
box 0 0 1 1
use contact_7  contact_7_523
timestamp 1624857261
transform 1 0 6466 0 1 14959
box 0 0 1 1
use contact_19  contact_19_521
timestamp 1624857261
transform 1 0 6899 0 1 14964
box 0 0 1 1
use contact_7  contact_7_521
timestamp 1624857261
transform 1 0 6898 0 1 14959
box 0 0 1 1
use contact_19  contact_19_178
timestamp 1624857261
transform 1 0 7281 0 1 14978
box 0 0 1 1
use contact_7  contact_7_178
timestamp 1624857261
transform 1 0 7280 0 1 14973
box 0 0 1 1
use contact_17  contact_17_269
timestamp 1624857261
transform 1 0 4664 0 1 15062
box 0 0 1 1
use contact_17  contact_17_268
timestamp 1624857261
transform 1 0 4904 0 1 15174
box 0 0 1 1
use contact_17  contact_17_267
timestamp 1624857261
transform 1 0 5304 0 1 15264
box 0 0 1 1
use contact_19  contact_19_179
timestamp 1624857261
transform 1 0 6042 0 1 15022
box 0 0 1 1
use contact_7  contact_7_179
timestamp 1624857261
transform 1 0 6041 0 1 15017
box 0 0 1 1
use and3_dec  and3_dec_89
timestamp 1624857261
transform 1 0 5803 0 1 15010
box 0 -60 2072 490
use contact_17  contact_17_264
timestamp 1624857261
transform 1 0 5304 0 1 15488
box 0 0 1 1
use contact_19  contact_19_520
timestamp 1624857261
transform 1 0 6467 0 1 15396
box 0 0 1 1
use contact_7  contact_7_520
timestamp 1624857261
transform 1 0 6466 0 1 15391
box 0 0 1 1
use contact_19  contact_19_518
timestamp 1624857261
transform 1 0 6899 0 1 15396
box 0 0 1 1
use contact_7  contact_7_518
timestamp 1624857261
transform 1 0 6898 0 1 15391
box 0 0 1 1
use contact_19  contact_19_177
timestamp 1624857261
transform 1 0 6042 0 1 15396
box 0 0 1 1
use contact_7  contact_7_177
timestamp 1624857261
transform 1 0 6041 0 1 15391
box 0 0 1 1
use contact_19  contact_19_176
timestamp 1624857261
transform 1 0 7281 0 1 15373
box 0 0 1 1
use contact_7  contact_7_176
timestamp 1624857261
transform 1 0 7280 0 1 15368
box 0 0 1 1
use contact_17  contact_17_265
timestamp 1624857261
transform 1 0 4904 0 1 15578
box 0 0 1 1
use contact_17  contact_17_266
timestamp 1624857261
transform 1 0 4744 0 1 15690
box 0 0 1 1
use contact_7  contact_7_175
timestamp 1624857261
transform 1 0 6041 0 1 15807
box 0 0 1 1
use contact_19  contact_19_175
timestamp 1624857261
transform 1 0 6042 0 1 15812
box 0 0 1 1
use contact_7  contact_7_517
timestamp 1624857261
transform 1 0 6466 0 1 15749
box 0 0 1 1
use contact_19  contact_19_517
timestamp 1624857261
transform 1 0 6467 0 1 15754
box 0 0 1 1
use contact_7  contact_7_515
timestamp 1624857261
transform 1 0 6898 0 1 15749
box 0 0 1 1
use contact_19  contact_19_515
timestamp 1624857261
transform 1 0 6899 0 1 15754
box 0 0 1 1
use contact_7  contact_7_174
timestamp 1624857261
transform 1 0 7280 0 1 15763
box 0 0 1 1
use contact_19  contact_19_174
timestamp 1624857261
transform 1 0 7281 0 1 15768
box 0 0 1 1
use and3_dec  and3_dec_88
timestamp 1624857261
transform 1 0 5803 0 -1 15800
box 0 -60 2072 490
use and3_dec  and3_dec_87
timestamp 1624857261
transform 1 0 5803 0 1 15800
box 0 -60 2072 490
use contact_17  contact_17_263
timestamp 1624857261
transform 1 0 4504 0 1 15852
box 0 0 1 1
use contact_17  contact_17_262
timestamp 1624857261
transform 1 0 4984 0 1 15964
box 0 0 1 1
use contact_17  contact_17_261
timestamp 1624857261
transform 1 0 5304 0 1 16054
box 0 0 1 1
use contact_17  contact_17_258
timestamp 1624857261
transform 1 0 5304 0 1 16278
box 0 0 1 1
use contact_19  contact_19_514
timestamp 1624857261
transform 1 0 6467 0 1 16186
box 0 0 1 1
use contact_7  contact_7_514
timestamp 1624857261
transform 1 0 6466 0 1 16181
box 0 0 1 1
use contact_19  contact_19_512
timestamp 1624857261
transform 1 0 6899 0 1 16186
box 0 0 1 1
use contact_7  contact_7_512
timestamp 1624857261
transform 1 0 6898 0 1 16181
box 0 0 1 1
use contact_19  contact_19_173
timestamp 1624857261
transform 1 0 6042 0 1 16186
box 0 0 1 1
use contact_7  contact_7_173
timestamp 1624857261
transform 1 0 6041 0 1 16181
box 0 0 1 1
use contact_19  contact_19_172
timestamp 1624857261
transform 1 0 7281 0 1 16163
box 0 0 1 1
use contact_7  contact_7_172
timestamp 1624857261
transform 1 0 7280 0 1 16158
box 0 0 1 1
use and3_dec  and3_dec_86
timestamp 1624857261
transform 1 0 5803 0 -1 16590
box 0 -60 2072 490
use contact_7  contact_7_531
timestamp 1624857261
transform 1 0 7676 0 1 13788
box 0 0 1 1
use contact_19  contact_19_531
timestamp 1624857261
transform 1 0 7677 0 1 13793
box 0 0 1 1
use contact_7  contact_7_534
timestamp 1624857261
transform 1 0 7676 0 1 13393
box 0 0 1 1
use contact_19  contact_19_534
timestamp 1624857261
transform 1 0 7677 0 1 13398
box 0 0 1 1
use contact_7  contact_7_525
timestamp 1624857261
transform 1 0 7676 0 1 14578
box 0 0 1 1
use contact_19  contact_19_525
timestamp 1624857261
transform 1 0 7677 0 1 14583
box 0 0 1 1
use contact_7  contact_7_528
timestamp 1624857261
transform 1 0 7676 0 1 14183
box 0 0 1 1
use contact_19  contact_19_528
timestamp 1624857261
transform 1 0 7677 0 1 14188
box 0 0 1 1
use contact_7  contact_7_519
timestamp 1624857261
transform 1 0 7676 0 1 15368
box 0 0 1 1
use contact_19  contact_19_519
timestamp 1624857261
transform 1 0 7677 0 1 15373
box 0 0 1 1
use contact_7  contact_7_522
timestamp 1624857261
transform 1 0 7676 0 1 14973
box 0 0 1 1
use contact_19  contact_19_522
timestamp 1624857261
transform 1 0 7677 0 1 14978
box 0 0 1 1
use contact_7  contact_7_513
timestamp 1624857261
transform 1 0 7676 0 1 16158
box 0 0 1 1
use contact_19  contact_19_513
timestamp 1624857261
transform 1 0 7677 0 1 16163
box 0 0 1 1
use contact_7  contact_7_516
timestamp 1624857261
transform 1 0 7676 0 1 15763
box 0 0 1 1
use contact_19  contact_19_516
timestamp 1624857261
transform 1 0 7677 0 1 15768
box 0 0 1 1
use contact_17  contact_17_260
timestamp 1624857261
transform 1 0 4584 0 1 16480
box 0 0 1 1
use contact_17  contact_17_259
timestamp 1624857261
transform 1 0 4984 0 1 16368
box 0 0 1 1
use contact_7  contact_7_171
timestamp 1624857261
transform 1 0 6041 0 1 16597
box 0 0 1 1
use contact_19  contact_19_171
timestamp 1624857261
transform 1 0 6042 0 1 16602
box 0 0 1 1
use contact_7  contact_7_511
timestamp 1624857261
transform 1 0 6466 0 1 16539
box 0 0 1 1
use contact_19  contact_19_511
timestamp 1624857261
transform 1 0 6467 0 1 16544
box 0 0 1 1
use contact_7  contact_7_509
timestamp 1624857261
transform 1 0 6898 0 1 16539
box 0 0 1 1
use contact_19  contact_19_509
timestamp 1624857261
transform 1 0 6899 0 1 16544
box 0 0 1 1
use contact_7  contact_7_170
timestamp 1624857261
transform 1 0 7280 0 1 16553
box 0 0 1 1
use contact_19  contact_19_170
timestamp 1624857261
transform 1 0 7281 0 1 16558
box 0 0 1 1
use contact_17  contact_17_257
timestamp 1624857261
transform 1 0 4664 0 1 16642
box 0 0 1 1
use contact_17  contact_17_256
timestamp 1624857261
transform 1 0 4984 0 1 16754
box 0 0 1 1
use contact_17  contact_17_255
timestamp 1624857261
transform 1 0 5304 0 1 16844
box 0 0 1 1
use and3_dec  and3_dec_85
timestamp 1624857261
transform 1 0 5803 0 1 16590
box 0 -60 2072 490
use and3_dec  and3_dec_84
timestamp 1624857261
transform 1 0 5803 0 -1 17380
box 0 -60 2072 490
use contact_17  contact_17_252
timestamp 1624857261
transform 1 0 5304 0 1 17068
box 0 0 1 1
use contact_17  contact_17_253
timestamp 1624857261
transform 1 0 4984 0 1 17158
box 0 0 1 1
use contact_7  contact_7_169
timestamp 1624857261
transform 1 0 6041 0 1 16971
box 0 0 1 1
use contact_19  contact_19_169
timestamp 1624857261
transform 1 0 6042 0 1 16976
box 0 0 1 1
use contact_7  contact_7_508
timestamp 1624857261
transform 1 0 6466 0 1 16971
box 0 0 1 1
use contact_19  contact_19_508
timestamp 1624857261
transform 1 0 6467 0 1 16976
box 0 0 1 1
use contact_7  contact_7_506
timestamp 1624857261
transform 1 0 6898 0 1 16971
box 0 0 1 1
use contact_19  contact_19_506
timestamp 1624857261
transform 1 0 6899 0 1 16976
box 0 0 1 1
use contact_7  contact_7_168
timestamp 1624857261
transform 1 0 7280 0 1 16948
box 0 0 1 1
use contact_19  contact_19_168
timestamp 1624857261
transform 1 0 7281 0 1 16953
box 0 0 1 1
use contact_17  contact_17_251
timestamp 1624857261
transform 1 0 4504 0 1 17432
box 0 0 1 1
use contact_17  contact_17_254
timestamp 1624857261
transform 1 0 4744 0 1 17270
box 0 0 1 1
use contact_7  contact_7_167
timestamp 1624857261
transform 1 0 6041 0 1 17387
box 0 0 1 1
use contact_19  contact_19_167
timestamp 1624857261
transform 1 0 6042 0 1 17392
box 0 0 1 1
use contact_7  contact_7_505
timestamp 1624857261
transform 1 0 6466 0 1 17329
box 0 0 1 1
use contact_19  contact_19_505
timestamp 1624857261
transform 1 0 6467 0 1 17334
box 0 0 1 1
use contact_7  contact_7_503
timestamp 1624857261
transform 1 0 6898 0 1 17329
box 0 0 1 1
use contact_19  contact_19_503
timestamp 1624857261
transform 1 0 6899 0 1 17334
box 0 0 1 1
use contact_7  contact_7_166
timestamp 1624857261
transform 1 0 7280 0 1 17343
box 0 0 1 1
use contact_19  contact_19_166
timestamp 1624857261
transform 1 0 7281 0 1 17348
box 0 0 1 1
use and3_dec  and3_dec_83
timestamp 1624857261
transform 1 0 5803 0 1 17380
box 0 -60 2072 490
use contact_17  contact_17_250
timestamp 1624857261
transform 1 0 5064 0 1 17544
box 0 0 1 1
use contact_17  contact_17_249
timestamp 1624857261
transform 1 0 5304 0 1 17634
box 0 0 1 1
use contact_17  contact_17_246
timestamp 1624857261
transform 1 0 5304 0 1 17858
box 0 0 1 1
use contact_17  contact_17_247
timestamp 1624857261
transform 1 0 5064 0 1 17948
box 0 0 1 1
use contact_7  contact_7_165
timestamp 1624857261
transform 1 0 6041 0 1 17761
box 0 0 1 1
use contact_19  contact_19_165
timestamp 1624857261
transform 1 0 6042 0 1 17766
box 0 0 1 1
use contact_7  contact_7_502
timestamp 1624857261
transform 1 0 6466 0 1 17761
box 0 0 1 1
use contact_19  contact_19_502
timestamp 1624857261
transform 1 0 6467 0 1 17766
box 0 0 1 1
use contact_7  contact_7_500
timestamp 1624857261
transform 1 0 6898 0 1 17761
box 0 0 1 1
use contact_19  contact_19_500
timestamp 1624857261
transform 1 0 6899 0 1 17766
box 0 0 1 1
use contact_7  contact_7_164
timestamp 1624857261
transform 1 0 7280 0 1 17738
box 0 0 1 1
use contact_19  contact_19_164
timestamp 1624857261
transform 1 0 7281 0 1 17743
box 0 0 1 1
use and3_dec  and3_dec_82
timestamp 1624857261
transform 1 0 5803 0 -1 18170
box 0 -60 2072 490
use contact_17  contact_17_245
timestamp 1624857261
transform 1 0 4664 0 1 18222
box 0 0 1 1
use contact_17  contact_17_248
timestamp 1624857261
transform 1 0 4584 0 1 18060
box 0 0 1 1
use contact_7  contact_7_163
timestamp 1624857261
transform 1 0 6041 0 1 18177
box 0 0 1 1
use contact_19  contact_19_163
timestamp 1624857261
transform 1 0 6042 0 1 18182
box 0 0 1 1
use contact_7  contact_7_499
timestamp 1624857261
transform 1 0 6466 0 1 18119
box 0 0 1 1
use contact_19  contact_19_499
timestamp 1624857261
transform 1 0 6467 0 1 18124
box 0 0 1 1
use contact_7  contact_7_497
timestamp 1624857261
transform 1 0 6898 0 1 18119
box 0 0 1 1
use contact_19  contact_19_497
timestamp 1624857261
transform 1 0 6899 0 1 18124
box 0 0 1 1
use contact_7  contact_7_162
timestamp 1624857261
transform 1 0 7280 0 1 18133
box 0 0 1 1
use contact_19  contact_19_162
timestamp 1624857261
transform 1 0 7281 0 1 18138
box 0 0 1 1
use contact_17  contact_17_244
timestamp 1624857261
transform 1 0 5064 0 1 18334
box 0 0 1 1
use contact_17  contact_17_243
timestamp 1624857261
transform 1 0 5304 0 1 18424
box 0 0 1 1
use contact_19  contact_19_160
timestamp 1624857261
transform 1 0 7281 0 1 18533
box 0 0 1 1
use contact_7  contact_7_160
timestamp 1624857261
transform 1 0 7280 0 1 18528
box 0 0 1 1
use and3_dec  and3_dec_81
timestamp 1624857261
transform 1 0 5803 0 1 18170
box 0 -60 2072 490
use and3_dec  and3_dec_80
timestamp 1624857261
transform 1 0 5803 0 -1 18960
box 0 -60 2072 490
use contact_17  contact_17_241
timestamp 1624857261
transform 1 0 5064 0 1 18738
box 0 0 1 1
use contact_17  contact_17_240
timestamp 1624857261
transform 1 0 5304 0 1 18648
box 0 0 1 1
use contact_19  contact_19_496
timestamp 1624857261
transform 1 0 6467 0 1 18556
box 0 0 1 1
use contact_7  contact_7_496
timestamp 1624857261
transform 1 0 6466 0 1 18551
box 0 0 1 1
use contact_19  contact_19_494
timestamp 1624857261
transform 1 0 6899 0 1 18556
box 0 0 1 1
use contact_7  contact_7_494
timestamp 1624857261
transform 1 0 6898 0 1 18551
box 0 0 1 1
use contact_19  contact_19_161
timestamp 1624857261
transform 1 0 6042 0 1 18556
box 0 0 1 1
use contact_7  contact_7_161
timestamp 1624857261
transform 1 0 6041 0 1 18551
box 0 0 1 1
use contact_17  contact_17_239
timestamp 1624857261
transform 1 0 4504 0 1 19012
box 0 0 1 1
use contact_17  contact_17_242
timestamp 1624857261
transform 1 0 4744 0 1 18850
box 0 0 1 1
use contact_7  contact_7_159
timestamp 1624857261
transform 1 0 6041 0 1 18967
box 0 0 1 1
use contact_19  contact_19_159
timestamp 1624857261
transform 1 0 6042 0 1 18972
box 0 0 1 1
use contact_7  contact_7_493
timestamp 1624857261
transform 1 0 6466 0 1 18909
box 0 0 1 1
use contact_19  contact_19_493
timestamp 1624857261
transform 1 0 6467 0 1 18914
box 0 0 1 1
use contact_7  contact_7_491
timestamp 1624857261
transform 1 0 6898 0 1 18909
box 0 0 1 1
use contact_19  contact_19_491
timestamp 1624857261
transform 1 0 6899 0 1 18914
box 0 0 1 1
use contact_7  contact_7_158
timestamp 1624857261
transform 1 0 7280 0 1 18923
box 0 0 1 1
use contact_19  contact_19_158
timestamp 1624857261
transform 1 0 7281 0 1 18928
box 0 0 1 1
use and3_dec  and3_dec_79
timestamp 1624857261
transform 1 0 5803 0 1 18960
box 0 -60 2072 490
use contact_17  contact_17_238
timestamp 1624857261
transform 1 0 4824 0 1 19124
box 0 0 1 1
use contact_17  contact_17_237
timestamp 1624857261
transform 1 0 5384 0 1 19214
box 0 0 1 1
use contact_7  contact_7_157
timestamp 1624857261
transform 1 0 6041 0 1 19341
box 0 0 1 1
use contact_19  contact_19_157
timestamp 1624857261
transform 1 0 6042 0 1 19346
box 0 0 1 1
use contact_7  contact_7_490
timestamp 1624857261
transform 1 0 6466 0 1 19341
box 0 0 1 1
use contact_19  contact_19_490
timestamp 1624857261
transform 1 0 6467 0 1 19346
box 0 0 1 1
use contact_7  contact_7_488
timestamp 1624857261
transform 1 0 6898 0 1 19341
box 0 0 1 1
use contact_19  contact_19_488
timestamp 1624857261
transform 1 0 6899 0 1 19346
box 0 0 1 1
use contact_7  contact_7_156
timestamp 1624857261
transform 1 0 7280 0 1 19318
box 0 0 1 1
use contact_19  contact_19_156
timestamp 1624857261
transform 1 0 7281 0 1 19323
box 0 0 1 1
use contact_17  contact_17_235
timestamp 1624857261
transform 1 0 4824 0 1 19528
box 0 0 1 1
use contact_17  contact_17_234
timestamp 1624857261
transform 1 0 5384 0 1 19438
box 0 0 1 1
use and3_dec  and3_dec_78
timestamp 1624857261
transform 1 0 5803 0 -1 19750
box 0 -60 2072 490
use contact_7  contact_7_507
timestamp 1624857261
transform 1 0 7676 0 1 16948
box 0 0 1 1
use contact_19  contact_19_507
timestamp 1624857261
transform 1 0 7677 0 1 16953
box 0 0 1 1
use contact_7  contact_7_510
timestamp 1624857261
transform 1 0 7676 0 1 16553
box 0 0 1 1
use contact_19  contact_19_510
timestamp 1624857261
transform 1 0 7677 0 1 16558
box 0 0 1 1
use contact_7  contact_7_501
timestamp 1624857261
transform 1 0 7676 0 1 17738
box 0 0 1 1
use contact_19  contact_19_501
timestamp 1624857261
transform 1 0 7677 0 1 17743
box 0 0 1 1
use contact_7  contact_7_504
timestamp 1624857261
transform 1 0 7676 0 1 17343
box 0 0 1 1
use contact_19  contact_19_504
timestamp 1624857261
transform 1 0 7677 0 1 17348
box 0 0 1 1
use contact_7  contact_7_492
timestamp 1624857261
transform 1 0 7676 0 1 18923
box 0 0 1 1
use contact_19  contact_19_492
timestamp 1624857261
transform 1 0 7677 0 1 18928
box 0 0 1 1
use contact_7  contact_7_495
timestamp 1624857261
transform 1 0 7676 0 1 18528
box 0 0 1 1
use contact_19  contact_19_495
timestamp 1624857261
transform 1 0 7677 0 1 18533
box 0 0 1 1
use contact_7  contact_7_498
timestamp 1624857261
transform 1 0 7676 0 1 18133
box 0 0 1 1
use contact_19  contact_19_498
timestamp 1624857261
transform 1 0 7677 0 1 18138
box 0 0 1 1
use contact_7  contact_7_489
timestamp 1624857261
transform 1 0 7676 0 1 19318
box 0 0 1 1
use contact_19  contact_19_489
timestamp 1624857261
transform 1 0 7677 0 1 19323
box 0 0 1 1
use contact_17  contact_17_233
timestamp 1624857261
transform 1 0 4664 0 1 19802
box 0 0 1 1
use contact_17  contact_17_236
timestamp 1624857261
transform 1 0 4584 0 1 19640
box 0 0 1 1
use contact_7  contact_7_155
timestamp 1624857261
transform 1 0 6041 0 1 19757
box 0 0 1 1
use contact_19  contact_19_155
timestamp 1624857261
transform 1 0 6042 0 1 19762
box 0 0 1 1
use contact_7  contact_7_487
timestamp 1624857261
transform 1 0 6466 0 1 19699
box 0 0 1 1
use contact_19  contact_19_487
timestamp 1624857261
transform 1 0 6467 0 1 19704
box 0 0 1 1
use contact_7  contact_7_485
timestamp 1624857261
transform 1 0 6898 0 1 19699
box 0 0 1 1
use contact_19  contact_19_485
timestamp 1624857261
transform 1 0 6899 0 1 19704
box 0 0 1 1
use contact_7  contact_7_154
timestamp 1624857261
transform 1 0 7280 0 1 19713
box 0 0 1 1
use contact_19  contact_19_154
timestamp 1624857261
transform 1 0 7281 0 1 19718
box 0 0 1 1
use contact_17  contact_17_232
timestamp 1624857261
transform 1 0 4824 0 1 19914
box 0 0 1 1
use contact_17  contact_17_231
timestamp 1624857261
transform 1 0 5384 0 1 20004
box 0 0 1 1
use contact_7  contact_7_153
timestamp 1624857261
transform 1 0 6041 0 1 20131
box 0 0 1 1
use contact_19  contact_19_153
timestamp 1624857261
transform 1 0 6042 0 1 20136
box 0 0 1 1
use contact_7  contact_7_484
timestamp 1624857261
transform 1 0 6466 0 1 20131
box 0 0 1 1
use contact_19  contact_19_484
timestamp 1624857261
transform 1 0 6467 0 1 20136
box 0 0 1 1
use contact_7  contact_7_482
timestamp 1624857261
transform 1 0 6898 0 1 20131
box 0 0 1 1
use contact_19  contact_19_482
timestamp 1624857261
transform 1 0 6899 0 1 20136
box 0 0 1 1
use contact_7  contact_7_152
timestamp 1624857261
transform 1 0 7280 0 1 20108
box 0 0 1 1
use contact_19  contact_19_152
timestamp 1624857261
transform 1 0 7281 0 1 20113
box 0 0 1 1
use and3_dec  and3_dec_77
timestamp 1624857261
transform 1 0 5803 0 1 19750
box 0 -60 2072 490
use and3_dec  and3_dec_76
timestamp 1624857261
transform 1 0 5803 0 -1 20540
box 0 -60 2072 490
use contact_17  contact_17_230
timestamp 1624857261
transform 1 0 4744 0 1 20430
box 0 0 1 1
use contact_17  contact_17_229
timestamp 1624857261
transform 1 0 4824 0 1 20318
box 0 0 1 1
use contact_17  contact_17_228
timestamp 1624857261
transform 1 0 5384 0 1 20228
box 0 0 1 1
use contact_17  contact_17_227
timestamp 1624857261
transform 1 0 4504 0 1 20592
box 0 0 1 1
use contact_17  contact_17_226
timestamp 1624857261
transform 1 0 4904 0 1 20704
box 0 0 1 1
use contact_7  contact_7_151
timestamp 1624857261
transform 1 0 6041 0 1 20547
box 0 0 1 1
use contact_19  contact_19_151
timestamp 1624857261
transform 1 0 6042 0 1 20552
box 0 0 1 1
use contact_7  contact_7_481
timestamp 1624857261
transform 1 0 6466 0 1 20489
box 0 0 1 1
use contact_19  contact_19_481
timestamp 1624857261
transform 1 0 6467 0 1 20494
box 0 0 1 1
use contact_7  contact_7_479
timestamp 1624857261
transform 1 0 6898 0 1 20489
box 0 0 1 1
use contact_19  contact_19_479
timestamp 1624857261
transform 1 0 6899 0 1 20494
box 0 0 1 1
use contact_7  contact_7_150
timestamp 1624857261
transform 1 0 7280 0 1 20503
box 0 0 1 1
use contact_19  contact_19_150
timestamp 1624857261
transform 1 0 7281 0 1 20508
box 0 0 1 1
use and3_dec  and3_dec_75
timestamp 1624857261
transform 1 0 5803 0 1 20540
box 0 -60 2072 490
use contact_17  contact_17_225
timestamp 1624857261
transform 1 0 5384 0 1 20794
box 0 0 1 1
use contact_19  contact_19_478
timestamp 1624857261
transform 1 0 6467 0 1 20926
box 0 0 1 1
use contact_7  contact_7_478
timestamp 1624857261
transform 1 0 6466 0 1 20921
box 0 0 1 1
use contact_19  contact_19_476
timestamp 1624857261
transform 1 0 6899 0 1 20926
box 0 0 1 1
use contact_7  contact_7_476
timestamp 1624857261
transform 1 0 6898 0 1 20921
box 0 0 1 1
use contact_19  contact_19_149
timestamp 1624857261
transform 1 0 6042 0 1 20926
box 0 0 1 1
use contact_7  contact_7_149
timestamp 1624857261
transform 1 0 6041 0 1 20921
box 0 0 1 1
use contact_19  contact_19_148
timestamp 1624857261
transform 1 0 7281 0 1 20903
box 0 0 1 1
use contact_7  contact_7_148
timestamp 1624857261
transform 1 0 7280 0 1 20898
box 0 0 1 1
use contact_17  contact_17_224
timestamp 1624857261
transform 1 0 4584 0 1 21220
box 0 0 1 1
use contact_17  contact_17_223
timestamp 1624857261
transform 1 0 4904 0 1 21108
box 0 0 1 1
use contact_17  contact_17_222
timestamp 1624857261
transform 1 0 5384 0 1 21018
box 0 0 1 1
use and3_dec  and3_dec_74
timestamp 1624857261
transform 1 0 5803 0 -1 21330
box 0 -60 2072 490
use and3_dec  and3_dec_73
timestamp 1624857261
transform 1 0 5803 0 1 21330
box 0 -60 2072 490
use contact_17  contact_17_220
timestamp 1624857261
transform 1 0 4904 0 1 21494
box 0 0 1 1
use contact_17  contact_17_221
timestamp 1624857261
transform 1 0 4664 0 1 21382
box 0 0 1 1
use contact_7  contact_7_147
timestamp 1624857261
transform 1 0 6041 0 1 21337
box 0 0 1 1
use contact_19  contact_19_147
timestamp 1624857261
transform 1 0 6042 0 1 21342
box 0 0 1 1
use contact_7  contact_7_475
timestamp 1624857261
transform 1 0 6466 0 1 21279
box 0 0 1 1
use contact_19  contact_19_475
timestamp 1624857261
transform 1 0 6467 0 1 21284
box 0 0 1 1
use contact_7  contact_7_473
timestamp 1624857261
transform 1 0 6898 0 1 21279
box 0 0 1 1
use contact_19  contact_19_473
timestamp 1624857261
transform 1 0 6899 0 1 21284
box 0 0 1 1
use contact_7  contact_7_146
timestamp 1624857261
transform 1 0 7280 0 1 21293
box 0 0 1 1
use contact_19  contact_19_146
timestamp 1624857261
transform 1 0 7281 0 1 21298
box 0 0 1 1
use contact_17  contact_17_216
timestamp 1624857261
transform 1 0 5384 0 1 21808
box 0 0 1 1
use contact_17  contact_17_219
timestamp 1624857261
transform 1 0 5384 0 1 21584
box 0 0 1 1
use contact_7  contact_7_145
timestamp 1624857261
transform 1 0 6041 0 1 21711
box 0 0 1 1
use contact_19  contact_19_145
timestamp 1624857261
transform 1 0 6042 0 1 21716
box 0 0 1 1
use contact_7  contact_7_472
timestamp 1624857261
transform 1 0 6466 0 1 21711
box 0 0 1 1
use contact_19  contact_19_472
timestamp 1624857261
transform 1 0 6467 0 1 21716
box 0 0 1 1
use contact_7  contact_7_470
timestamp 1624857261
transform 1 0 6898 0 1 21711
box 0 0 1 1
use contact_19  contact_19_470
timestamp 1624857261
transform 1 0 6899 0 1 21716
box 0 0 1 1
use contact_7  contact_7_144
timestamp 1624857261
transform 1 0 7280 0 1 21688
box 0 0 1 1
use contact_19  contact_19_144
timestamp 1624857261
transform 1 0 7281 0 1 21693
box 0 0 1 1
use and3_dec  and3_dec_72
timestamp 1624857261
transform 1 0 5803 0 -1 22120
box 0 -60 2072 490
use contact_17  contact_17_218
timestamp 1624857261
transform 1 0 4744 0 1 22010
box 0 0 1 1
use contact_17  contact_17_217
timestamp 1624857261
transform 1 0 4904 0 1 21898
box 0 0 1 1
use contact_19  contact_19_469
timestamp 1624857261
transform 1 0 6467 0 1 22074
box 0 0 1 1
use contact_7  contact_7_469
timestamp 1624857261
transform 1 0 6466 0 1 22069
box 0 0 1 1
use contact_19  contact_19_467
timestamp 1624857261
transform 1 0 6899 0 1 22074
box 0 0 1 1
use contact_7  contact_7_467
timestamp 1624857261
transform 1 0 6898 0 1 22069
box 0 0 1 1
use contact_19  contact_19_142
timestamp 1624857261
transform 1 0 7281 0 1 22088
box 0 0 1 1
use contact_7  contact_7_142
timestamp 1624857261
transform 1 0 7280 0 1 22083
box 0 0 1 1
use contact_17  contact_17_215
timestamp 1624857261
transform 1 0 4504 0 1 22172
box 0 0 1 1
use contact_17  contact_17_214
timestamp 1624857261
transform 1 0 4984 0 1 22284
box 0 0 1 1
use contact_17  contact_17_213
timestamp 1624857261
transform 1 0 5384 0 1 22374
box 0 0 1 1
use contact_19  contact_19_143
timestamp 1624857261
transform 1 0 6042 0 1 22132
box 0 0 1 1
use contact_7  contact_7_143
timestamp 1624857261
transform 1 0 6041 0 1 22127
box 0 0 1 1
use and3_dec  and3_dec_71
timestamp 1624857261
transform 1 0 5803 0 1 22120
box 0 -60 2072 490
use contact_17  contact_17_210
timestamp 1624857261
transform 1 0 5384 0 1 22598
box 0 0 1 1
use contact_19  contact_19_466
timestamp 1624857261
transform 1 0 6467 0 1 22506
box 0 0 1 1
use contact_7  contact_7_466
timestamp 1624857261
transform 1 0 6466 0 1 22501
box 0 0 1 1
use contact_19  contact_19_464
timestamp 1624857261
transform 1 0 6899 0 1 22506
box 0 0 1 1
use contact_7  contact_7_464
timestamp 1624857261
transform 1 0 6898 0 1 22501
box 0 0 1 1
use contact_19  contact_19_141
timestamp 1624857261
transform 1 0 6042 0 1 22506
box 0 0 1 1
use contact_7  contact_7_141
timestamp 1624857261
transform 1 0 6041 0 1 22501
box 0 0 1 1
use contact_19  contact_19_140
timestamp 1624857261
transform 1 0 7281 0 1 22483
box 0 0 1 1
use contact_7  contact_7_140
timestamp 1624857261
transform 1 0 7280 0 1 22478
box 0 0 1 1
use contact_17  contact_17_212
timestamp 1624857261
transform 1 0 4584 0 1 22800
box 0 0 1 1
use contact_17  contact_17_211
timestamp 1624857261
transform 1 0 4984 0 1 22688
box 0 0 1 1
use contact_19  contact_19_463
timestamp 1624857261
transform 1 0 6467 0 1 22864
box 0 0 1 1
use contact_7  contact_7_463
timestamp 1624857261
transform 1 0 6466 0 1 22859
box 0 0 1 1
use contact_19  contact_19_461
timestamp 1624857261
transform 1 0 6899 0 1 22864
box 0 0 1 1
use contact_7  contact_7_461
timestamp 1624857261
transform 1 0 6898 0 1 22859
box 0 0 1 1
use contact_19  contact_19_138
timestamp 1624857261
transform 1 0 7281 0 1 22878
box 0 0 1 1
use contact_7  contact_7_138
timestamp 1624857261
transform 1 0 7280 0 1 22873
box 0 0 1 1
use and3_dec  and3_dec_70
timestamp 1624857261
transform 1 0 5803 0 -1 22910
box 0 -60 2072 490
use and3_dec  and3_dec_69
timestamp 1624857261
transform 1 0 5803 0 1 22910
box 0 -60 2072 490
use contact_7  contact_7_483
timestamp 1624857261
transform 1 0 7676 0 1 20108
box 0 0 1 1
use contact_19  contact_19_483
timestamp 1624857261
transform 1 0 7677 0 1 20113
box 0 0 1 1
use contact_7  contact_7_486
timestamp 1624857261
transform 1 0 7676 0 1 19713
box 0 0 1 1
use contact_19  contact_19_486
timestamp 1624857261
transform 1 0 7677 0 1 19718
box 0 0 1 1
use contact_7  contact_7_477
timestamp 1624857261
transform 1 0 7676 0 1 20898
box 0 0 1 1
use contact_19  contact_19_477
timestamp 1624857261
transform 1 0 7677 0 1 20903
box 0 0 1 1
use contact_7  contact_7_480
timestamp 1624857261
transform 1 0 7676 0 1 20503
box 0 0 1 1
use contact_19  contact_19_480
timestamp 1624857261
transform 1 0 7677 0 1 20508
box 0 0 1 1
use contact_7  contact_7_468
timestamp 1624857261
transform 1 0 7676 0 1 22083
box 0 0 1 1
use contact_19  contact_19_468
timestamp 1624857261
transform 1 0 7677 0 1 22088
box 0 0 1 1
use contact_7  contact_7_471
timestamp 1624857261
transform 1 0 7676 0 1 21688
box 0 0 1 1
use contact_19  contact_19_471
timestamp 1624857261
transform 1 0 7677 0 1 21693
box 0 0 1 1
use contact_7  contact_7_474
timestamp 1624857261
transform 1 0 7676 0 1 21293
box 0 0 1 1
use contact_19  contact_19_474
timestamp 1624857261
transform 1 0 7677 0 1 21298
box 0 0 1 1
use contact_7  contact_7_462
timestamp 1624857261
transform 1 0 7676 0 1 22873
box 0 0 1 1
use contact_19  contact_19_462
timestamp 1624857261
transform 1 0 7677 0 1 22878
box 0 0 1 1
use contact_7  contact_7_465
timestamp 1624857261
transform 1 0 7676 0 1 22478
box 0 0 1 1
use contact_19  contact_19_465
timestamp 1624857261
transform 1 0 7677 0 1 22483
box 0 0 1 1
use contact_17  contact_17_209
timestamp 1624857261
transform 1 0 4664 0 1 22962
box 0 0 1 1
use contact_17  contact_17_208
timestamp 1624857261
transform 1 0 4984 0 1 23074
box 0 0 1 1
use contact_17  contact_17_207
timestamp 1624857261
transform 1 0 5384 0 1 23164
box 0 0 1 1
use contact_19  contact_19_139
timestamp 1624857261
transform 1 0 6042 0 1 22922
box 0 0 1 1
use contact_7  contact_7_139
timestamp 1624857261
transform 1 0 6041 0 1 22917
box 0 0 1 1
use contact_17  contact_17_204
timestamp 1624857261
transform 1 0 5384 0 1 23388
box 0 0 1 1
use contact_19  contact_19_460
timestamp 1624857261
transform 1 0 6467 0 1 23296
box 0 0 1 1
use contact_7  contact_7_460
timestamp 1624857261
transform 1 0 6466 0 1 23291
box 0 0 1 1
use contact_19  contact_19_458
timestamp 1624857261
transform 1 0 6899 0 1 23296
box 0 0 1 1
use contact_7  contact_7_458
timestamp 1624857261
transform 1 0 6898 0 1 23291
box 0 0 1 1
use contact_19  contact_19_137
timestamp 1624857261
transform 1 0 6042 0 1 23296
box 0 0 1 1
use contact_7  contact_7_137
timestamp 1624857261
transform 1 0 6041 0 1 23291
box 0 0 1 1
use contact_19  contact_19_136
timestamp 1624857261
transform 1 0 7281 0 1 23273
box 0 0 1 1
use contact_7  contact_7_136
timestamp 1624857261
transform 1 0 7280 0 1 23268
box 0 0 1 1
use and3_dec  and3_dec_68
timestamp 1624857261
transform 1 0 5803 0 -1 23700
box 0 -60 2072 490
use contact_17  contact_17_206
timestamp 1624857261
transform 1 0 4744 0 1 23590
box 0 0 1 1
use contact_17  contact_17_205
timestamp 1624857261
transform 1 0 4984 0 1 23478
box 0 0 1 1
use contact_7  contact_7_135
timestamp 1624857261
transform 1 0 6041 0 1 23707
box 0 0 1 1
use contact_19  contact_19_135
timestamp 1624857261
transform 1 0 6042 0 1 23712
box 0 0 1 1
use contact_7  contact_7_457
timestamp 1624857261
transform 1 0 6466 0 1 23649
box 0 0 1 1
use contact_19  contact_19_457
timestamp 1624857261
transform 1 0 6467 0 1 23654
box 0 0 1 1
use contact_7  contact_7_455
timestamp 1624857261
transform 1 0 6898 0 1 23649
box 0 0 1 1
use contact_19  contact_19_455
timestamp 1624857261
transform 1 0 6899 0 1 23654
box 0 0 1 1
use contact_7  contact_7_134
timestamp 1624857261
transform 1 0 7280 0 1 23663
box 0 0 1 1
use contact_19  contact_19_134
timestamp 1624857261
transform 1 0 7281 0 1 23668
box 0 0 1 1
use contact_17  contact_17_203
timestamp 1624857261
transform 1 0 4504 0 1 23752
box 0 0 1 1
use contact_17  contact_17_202
timestamp 1624857261
transform 1 0 5064 0 1 23864
box 0 0 1 1
use contact_17  contact_17_201
timestamp 1624857261
transform 1 0 5384 0 1 23954
box 0 0 1 1
use and3_dec  and3_dec_67
timestamp 1624857261
transform 1 0 5803 0 1 23700
box 0 -60 2072 490
use and3_dec  and3_dec_66
timestamp 1624857261
transform 1 0 5803 0 -1 24490
box 0 -60 2072 490
use contact_17  contact_17_199
timestamp 1624857261
transform 1 0 5064 0 1 24268
box 0 0 1 1
use contact_17  contact_17_198
timestamp 1624857261
transform 1 0 5384 0 1 24178
box 0 0 1 1
use contact_7  contact_7_133
timestamp 1624857261
transform 1 0 6041 0 1 24081
box 0 0 1 1
use contact_19  contact_19_133
timestamp 1624857261
transform 1 0 6042 0 1 24086
box 0 0 1 1
use contact_7  contact_7_454
timestamp 1624857261
transform 1 0 6466 0 1 24081
box 0 0 1 1
use contact_19  contact_19_454
timestamp 1624857261
transform 1 0 6467 0 1 24086
box 0 0 1 1
use contact_7  contact_7_452
timestamp 1624857261
transform 1 0 6898 0 1 24081
box 0 0 1 1
use contact_19  contact_19_452
timestamp 1624857261
transform 1 0 6899 0 1 24086
box 0 0 1 1
use contact_7  contact_7_132
timestamp 1624857261
transform 1 0 7280 0 1 24058
box 0 0 1 1
use contact_19  contact_19_132
timestamp 1624857261
transform 1 0 7281 0 1 24063
box 0 0 1 1
use contact_17  contact_17_197
timestamp 1624857261
transform 1 0 4664 0 1 24542
box 0 0 1 1
use contact_17  contact_17_200
timestamp 1624857261
transform 1 0 4584 0 1 24380
box 0 0 1 1
use contact_7  contact_7_131
timestamp 1624857261
transform 1 0 6041 0 1 24497
box 0 0 1 1
use contact_19  contact_19_131
timestamp 1624857261
transform 1 0 6042 0 1 24502
box 0 0 1 1
use contact_7  contact_7_451
timestamp 1624857261
transform 1 0 6466 0 1 24439
box 0 0 1 1
use contact_19  contact_19_451
timestamp 1624857261
transform 1 0 6467 0 1 24444
box 0 0 1 1
use contact_7  contact_7_449
timestamp 1624857261
transform 1 0 6898 0 1 24439
box 0 0 1 1
use contact_19  contact_19_449
timestamp 1624857261
transform 1 0 6899 0 1 24444
box 0 0 1 1
use contact_7  contact_7_130
timestamp 1624857261
transform 1 0 7280 0 1 24453
box 0 0 1 1
use contact_19  contact_19_130
timestamp 1624857261
transform 1 0 7281 0 1 24458
box 0 0 1 1
use and3_dec  and3_dec_65
timestamp 1624857261
transform 1 0 5803 0 1 24490
box 0 -60 2072 490
use contact_17  contact_17_196
timestamp 1624857261
transform 1 0 5064 0 1 24654
box 0 0 1 1
use contact_17  contact_17_195
timestamp 1624857261
transform 1 0 5384 0 1 24744
box 0 0 1 1
use contact_17  contact_17_193
timestamp 1624857261
transform 1 0 5064 0 1 25058
box 0 0 1 1
use contact_17  contact_17_192
timestamp 1624857261
transform 1 0 5384 0 1 24968
box 0 0 1 1
use contact_7  contact_7_129
timestamp 1624857261
transform 1 0 6041 0 1 24871
box 0 0 1 1
use contact_19  contact_19_129
timestamp 1624857261
transform 1 0 6042 0 1 24876
box 0 0 1 1
use contact_7  contact_7_448
timestamp 1624857261
transform 1 0 6466 0 1 24871
box 0 0 1 1
use contact_19  contact_19_448
timestamp 1624857261
transform 1 0 6467 0 1 24876
box 0 0 1 1
use contact_7  contact_7_446
timestamp 1624857261
transform 1 0 6898 0 1 24871
box 0 0 1 1
use contact_19  contact_19_446
timestamp 1624857261
transform 1 0 6899 0 1 24876
box 0 0 1 1
use contact_7  contact_7_128
timestamp 1624857261
transform 1 0 7280 0 1 24848
box 0 0 1 1
use contact_19  contact_19_128
timestamp 1624857261
transform 1 0 7281 0 1 24853
box 0 0 1 1
use and3_dec  and3_dec_64
timestamp 1624857261
transform 1 0 5803 0 -1 25280
box 0 -60 2072 490
use contact_17  contact_17_191
timestamp 1624857261
transform 1 0 4504 0 1 25332
box 0 0 1 1
use contact_17  contact_17_194
timestamp 1624857261
transform 1 0 4744 0 1 25170
box 0 0 1 1
use contact_7  contact_7_127
timestamp 1624857261
transform 1 0 6041 0 1 25287
box 0 0 1 1
use contact_19  contact_19_127
timestamp 1624857261
transform 1 0 6042 0 1 25292
box 0 0 1 1
use contact_7  contact_7_445
timestamp 1624857261
transform 1 0 6466 0 1 25229
box 0 0 1 1
use contact_19  contact_19_445
timestamp 1624857261
transform 1 0 6467 0 1 25234
box 0 0 1 1
use contact_7  contact_7_443
timestamp 1624857261
transform 1 0 6898 0 1 25229
box 0 0 1 1
use contact_19  contact_19_443
timestamp 1624857261
transform 1 0 6899 0 1 25234
box 0 0 1 1
use contact_7  contact_7_126
timestamp 1624857261
transform 1 0 7280 0 1 25243
box 0 0 1 1
use contact_19  contact_19_126
timestamp 1624857261
transform 1 0 7281 0 1 25248
box 0 0 1 1
use contact_17  contact_17_190
timestamp 1624857261
transform 1 0 4824 0 1 25444
box 0 0 1 1
use contact_17  contact_17_189
timestamp 1624857261
transform 1 0 5464 0 1 25534
box 0 0 1 1
use contact_7  contact_7_442
timestamp 1624857261
transform 1 0 6466 0 1 25661
box 0 0 1 1
use contact_7  contact_7_440
timestamp 1624857261
transform 1 0 6898 0 1 25661
box 0 0 1 1
use contact_7  contact_7_125
timestamp 1624857261
transform 1 0 6041 0 1 25661
box 0 0 1 1
use contact_19  contact_19_124
timestamp 1624857261
transform 1 0 7281 0 1 25643
box 0 0 1 1
use contact_7  contact_7_124
timestamp 1624857261
transform 1 0 7280 0 1 25638
box 0 0 1 1
use and3_dec  and3_dec_63
timestamp 1624857261
transform 1 0 5803 0 1 25280
box 0 -60 2072 490
use and3_dec  and3_dec_62
timestamp 1624857261
transform 1 0 5803 0 -1 26070
box 0 -60 2072 490
use contact_17  contact_17_187
timestamp 1624857261
transform 1 0 4824 0 1 25848
box 0 0 1 1
use contact_17  contact_17_186
timestamp 1624857261
transform 1 0 5464 0 1 25758
box 0 0 1 1
use contact_19  contact_19_442
timestamp 1624857261
transform 1 0 6467 0 1 25666
box 0 0 1 1
use contact_19  contact_19_440
timestamp 1624857261
transform 1 0 6899 0 1 25666
box 0 0 1 1
use contact_19  contact_19_125
timestamp 1624857261
transform 1 0 6042 0 1 25666
box 0 0 1 1
use contact_17  contact_17_185
timestamp 1624857261
transform 1 0 4664 0 1 26122
box 0 0 1 1
use contact_17  contact_17_188
timestamp 1624857261
transform 1 0 4584 0 1 25960
box 0 0 1 1
use contact_7  contact_7_123
timestamp 1624857261
transform 1 0 6041 0 1 26077
box 0 0 1 1
use contact_19  contact_19_123
timestamp 1624857261
transform 1 0 6042 0 1 26082
box 0 0 1 1
use contact_7  contact_7_439
timestamp 1624857261
transform 1 0 6466 0 1 26019
box 0 0 1 1
use contact_19  contact_19_439
timestamp 1624857261
transform 1 0 6467 0 1 26024
box 0 0 1 1
use contact_7  contact_7_437
timestamp 1624857261
transform 1 0 6898 0 1 26019
box 0 0 1 1
use contact_19  contact_19_437
timestamp 1624857261
transform 1 0 6899 0 1 26024
box 0 0 1 1
use contact_7  contact_7_122
timestamp 1624857261
transform 1 0 7280 0 1 26033
box 0 0 1 1
use contact_19  contact_19_122
timestamp 1624857261
transform 1 0 7281 0 1 26038
box 0 0 1 1
use and3_dec  and3_dec_61
timestamp 1624857261
transform 1 0 5803 0 1 26070
box 0 -60 2072 490
use contact_7  contact_7_456
timestamp 1624857261
transform 1 0 7676 0 1 23663
box 0 0 1 1
use contact_19  contact_19_456
timestamp 1624857261
transform 1 0 7677 0 1 23668
box 0 0 1 1
use contact_7  contact_7_459
timestamp 1624857261
transform 1 0 7676 0 1 23268
box 0 0 1 1
use contact_19  contact_19_459
timestamp 1624857261
transform 1 0 7677 0 1 23273
box 0 0 1 1
use contact_7  contact_7_450
timestamp 1624857261
transform 1 0 7676 0 1 24453
box 0 0 1 1
use contact_19  contact_19_450
timestamp 1624857261
transform 1 0 7677 0 1 24458
box 0 0 1 1
use contact_7  contact_7_453
timestamp 1624857261
transform 1 0 7676 0 1 24058
box 0 0 1 1
use contact_19  contact_19_453
timestamp 1624857261
transform 1 0 7677 0 1 24063
box 0 0 1 1
use contact_7  contact_7_444
timestamp 1624857261
transform 1 0 7676 0 1 25243
box 0 0 1 1
use contact_19  contact_19_444
timestamp 1624857261
transform 1 0 7677 0 1 25248
box 0 0 1 1
use contact_7  contact_7_447
timestamp 1624857261
transform 1 0 7676 0 1 24848
box 0 0 1 1
use contact_19  contact_19_447
timestamp 1624857261
transform 1 0 7677 0 1 24853
box 0 0 1 1
use contact_7  contact_7_438
timestamp 1624857261
transform 1 0 7676 0 1 26033
box 0 0 1 1
use contact_19  contact_19_438
timestamp 1624857261
transform 1 0 7677 0 1 26038
box 0 0 1 1
use contact_7  contact_7_441
timestamp 1624857261
transform 1 0 7676 0 1 25638
box 0 0 1 1
use contact_19  contact_19_441
timestamp 1624857261
transform 1 0 7677 0 1 25643
box 0 0 1 1
use contact_17  contact_17_184
timestamp 1624857261
transform 1 0 4824 0 1 26234
box 0 0 1 1
use contact_17  contact_17_183
timestamp 1624857261
transform 1 0 5464 0 1 26324
box 0 0 1 1
use contact_7  contact_7_121
timestamp 1624857261
transform 1 0 6041 0 1 26451
box 0 0 1 1
use contact_19  contact_19_121
timestamp 1624857261
transform 1 0 6042 0 1 26456
box 0 0 1 1
use contact_7  contact_7_436
timestamp 1624857261
transform 1 0 6466 0 1 26451
box 0 0 1 1
use contact_19  contact_19_436
timestamp 1624857261
transform 1 0 6467 0 1 26456
box 0 0 1 1
use contact_7  contact_7_434
timestamp 1624857261
transform 1 0 6898 0 1 26451
box 0 0 1 1
use contact_19  contact_19_434
timestamp 1624857261
transform 1 0 6899 0 1 26456
box 0 0 1 1
use contact_7  contact_7_120
timestamp 1624857261
transform 1 0 7280 0 1 26428
box 0 0 1 1
use contact_19  contact_19_120
timestamp 1624857261
transform 1 0 7281 0 1 26433
box 0 0 1 1
use contact_17  contact_17_181
timestamp 1624857261
transform 1 0 4824 0 1 26638
box 0 0 1 1
use contact_17  contact_17_180
timestamp 1624857261
transform 1 0 5464 0 1 26548
box 0 0 1 1
use and3_dec  and3_dec_60
timestamp 1624857261
transform 1 0 5803 0 -1 26860
box 0 -60 2072 490
use contact_17  contact_17_179
timestamp 1624857261
transform 1 0 4504 0 1 26912
box 0 0 1 1
use contact_17  contact_17_182
timestamp 1624857261
transform 1 0 4744 0 1 26750
box 0 0 1 1
use contact_7  contact_7_119
timestamp 1624857261
transform 1 0 6041 0 1 26867
box 0 0 1 1
use contact_19  contact_19_119
timestamp 1624857261
transform 1 0 6042 0 1 26872
box 0 0 1 1
use contact_7  contact_7_433
timestamp 1624857261
transform 1 0 6466 0 1 26809
box 0 0 1 1
use contact_19  contact_19_433
timestamp 1624857261
transform 1 0 6467 0 1 26814
box 0 0 1 1
use contact_7  contact_7_431
timestamp 1624857261
transform 1 0 6898 0 1 26809
box 0 0 1 1
use contact_19  contact_19_431
timestamp 1624857261
transform 1 0 6899 0 1 26814
box 0 0 1 1
use contact_7  contact_7_118
timestamp 1624857261
transform 1 0 7280 0 1 26823
box 0 0 1 1
use contact_19  contact_19_118
timestamp 1624857261
transform 1 0 7281 0 1 26828
box 0 0 1 1
use contact_17  contact_17_178
timestamp 1624857261
transform 1 0 4904 0 1 27024
box 0 0 1 1
use contact_17  contact_17_177
timestamp 1624857261
transform 1 0 5464 0 1 27114
box 0 0 1 1
use contact_7  contact_7_117
timestamp 1624857261
transform 1 0 6041 0 1 27241
box 0 0 1 1
use contact_19  contact_19_117
timestamp 1624857261
transform 1 0 6042 0 1 27246
box 0 0 1 1
use contact_7  contact_7_430
timestamp 1624857261
transform 1 0 6466 0 1 27241
box 0 0 1 1
use contact_19  contact_19_430
timestamp 1624857261
transform 1 0 6467 0 1 27246
box 0 0 1 1
use contact_7  contact_7_428
timestamp 1624857261
transform 1 0 6898 0 1 27241
box 0 0 1 1
use contact_19  contact_19_428
timestamp 1624857261
transform 1 0 6899 0 1 27246
box 0 0 1 1
use contact_7  contact_7_116
timestamp 1624857261
transform 1 0 7280 0 1 27218
box 0 0 1 1
use contact_19  contact_19_116
timestamp 1624857261
transform 1 0 7281 0 1 27223
box 0 0 1 1
use and3_dec  and3_dec_59
timestamp 1624857261
transform 1 0 5803 0 1 26860
box 0 -60 2072 490
use and3_dec  and3_dec_58
timestamp 1624857261
transform 1 0 5803 0 -1 27650
box 0 -60 2072 490
use contact_17  contact_17_176
timestamp 1624857261
transform 1 0 4584 0 1 27540
box 0 0 1 1
use contact_17  contact_17_175
timestamp 1624857261
transform 1 0 4904 0 1 27428
box 0 0 1 1
use contact_17  contact_17_174
timestamp 1624857261
transform 1 0 5464 0 1 27338
box 0 0 1 1
use contact_17  contact_17_172
timestamp 1624857261
transform 1 0 4904 0 1 27814
box 0 0 1 1
use contact_17  contact_17_173
timestamp 1624857261
transform 1 0 4664 0 1 27702
box 0 0 1 1
use contact_7  contact_7_115
timestamp 1624857261
transform 1 0 6041 0 1 27657
box 0 0 1 1
use contact_19  contact_19_115
timestamp 1624857261
transform 1 0 6042 0 1 27662
box 0 0 1 1
use contact_7  contact_7_427
timestamp 1624857261
transform 1 0 6466 0 1 27599
box 0 0 1 1
use contact_19  contact_19_427
timestamp 1624857261
transform 1 0 6467 0 1 27604
box 0 0 1 1
use contact_7  contact_7_425
timestamp 1624857261
transform 1 0 6898 0 1 27599
box 0 0 1 1
use contact_19  contact_19_425
timestamp 1624857261
transform 1 0 6899 0 1 27604
box 0 0 1 1
use contact_7  contact_7_114
timestamp 1624857261
transform 1 0 7280 0 1 27613
box 0 0 1 1
use contact_19  contact_19_114
timestamp 1624857261
transform 1 0 7281 0 1 27618
box 0 0 1 1
use and3_dec  and3_dec_57
timestamp 1624857261
transform 1 0 5803 0 1 27650
box 0 -60 2072 490
use contact_17  contact_17_171
timestamp 1624857261
transform 1 0 5464 0 1 27904
box 0 0 1 1
use contact_19  contact_19_424
timestamp 1624857261
transform 1 0 6467 0 1 28036
box 0 0 1 1
use contact_7  contact_7_424
timestamp 1624857261
transform 1 0 6466 0 1 28031
box 0 0 1 1
use contact_19  contact_19_422
timestamp 1624857261
transform 1 0 6899 0 1 28036
box 0 0 1 1
use contact_7  contact_7_422
timestamp 1624857261
transform 1 0 6898 0 1 28031
box 0 0 1 1
use contact_19  contact_19_113
timestamp 1624857261
transform 1 0 6042 0 1 28036
box 0 0 1 1
use contact_7  contact_7_113
timestamp 1624857261
transform 1 0 6041 0 1 28031
box 0 0 1 1
use contact_19  contact_19_112
timestamp 1624857261
transform 1 0 7281 0 1 28013
box 0 0 1 1
use contact_7  contact_7_112
timestamp 1624857261
transform 1 0 7280 0 1 28008
box 0 0 1 1
use contact_17  contact_17_170
timestamp 1624857261
transform 1 0 4744 0 1 28330
box 0 0 1 1
use contact_17  contact_17_169
timestamp 1624857261
transform 1 0 4904 0 1 28218
box 0 0 1 1
use contact_17  contact_17_168
timestamp 1624857261
transform 1 0 5464 0 1 28128
box 0 0 1 1
use contact_7  contact_7_421
timestamp 1624857261
transform 1 0 6466 0 1 28389
box 0 0 1 1
use contact_7  contact_7_419
timestamp 1624857261
transform 1 0 6898 0 1 28389
box 0 0 1 1
use and3_dec  and3_dec_56
timestamp 1624857261
transform 1 0 5803 0 -1 28440
box 0 -60 2072 490
use and3_dec  and3_dec_55
timestamp 1624857261
transform 1 0 5803 0 1 28440
box 0 -60 2072 490
use contact_17  contact_17_167
timestamp 1624857261
transform 1 0 4504 0 1 28492
box 0 0 1 1
use contact_17  contact_17_166
timestamp 1624857261
transform 1 0 4984 0 1 28604
box 0 0 1 1
use contact_19  contact_19_421
timestamp 1624857261
transform 1 0 6467 0 1 28394
box 0 0 1 1
use contact_19  contact_19_419
timestamp 1624857261
transform 1 0 6899 0 1 28394
box 0 0 1 1
use contact_19  contact_19_111
timestamp 1624857261
transform 1 0 6042 0 1 28452
box 0 0 1 1
use contact_7  contact_7_111
timestamp 1624857261
transform 1 0 6041 0 1 28447
box 0 0 1 1
use contact_19  contact_19_110
timestamp 1624857261
transform 1 0 7281 0 1 28408
box 0 0 1 1
use contact_7  contact_7_110
timestamp 1624857261
transform 1 0 7280 0 1 28403
box 0 0 1 1
use contact_17  contact_17_162
timestamp 1624857261
transform 1 0 5464 0 1 28918
box 0 0 1 1
use contact_17  contact_17_165
timestamp 1624857261
transform 1 0 5464 0 1 28694
box 0 0 1 1
use contact_7  contact_7_109
timestamp 1624857261
transform 1 0 6041 0 1 28821
box 0 0 1 1
use contact_19  contact_19_109
timestamp 1624857261
transform 1 0 6042 0 1 28826
box 0 0 1 1
use contact_7  contact_7_418
timestamp 1624857261
transform 1 0 6466 0 1 28821
box 0 0 1 1
use contact_19  contact_19_418
timestamp 1624857261
transform 1 0 6467 0 1 28826
box 0 0 1 1
use contact_7  contact_7_416
timestamp 1624857261
transform 1 0 6898 0 1 28821
box 0 0 1 1
use contact_19  contact_19_416
timestamp 1624857261
transform 1 0 6899 0 1 28826
box 0 0 1 1
use contact_7  contact_7_108
timestamp 1624857261
transform 1 0 7280 0 1 28798
box 0 0 1 1
use contact_19  contact_19_108
timestamp 1624857261
transform 1 0 7281 0 1 28803
box 0 0 1 1
use and3_dec  and3_dec_54
timestamp 1624857261
transform 1 0 5803 0 -1 29230
box 0 -60 2072 490
use contact_17  contact_17_164
timestamp 1624857261
transform 1 0 4584 0 1 29120
box 0 0 1 1
use contact_17  contact_17_163
timestamp 1624857261
transform 1 0 4984 0 1 29008
box 0 0 1 1
use contact_19  contact_19_415
timestamp 1624857261
transform 1 0 6467 0 1 29184
box 0 0 1 1
use contact_7  contact_7_415
timestamp 1624857261
transform 1 0 6466 0 1 29179
box 0 0 1 1
use contact_19  contact_19_413
timestamp 1624857261
transform 1 0 6899 0 1 29184
box 0 0 1 1
use contact_7  contact_7_413
timestamp 1624857261
transform 1 0 6898 0 1 29179
box 0 0 1 1
use contact_19  contact_19_106
timestamp 1624857261
transform 1 0 7281 0 1 29198
box 0 0 1 1
use contact_7  contact_7_106
timestamp 1624857261
transform 1 0 7280 0 1 29193
box 0 0 1 1
use contact_17  contact_17_161
timestamp 1624857261
transform 1 0 4664 0 1 29282
box 0 0 1 1
use contact_17  contact_17_160
timestamp 1624857261
transform 1 0 4984 0 1 29394
box 0 0 1 1
use contact_19  contact_19_107
timestamp 1624857261
transform 1 0 6042 0 1 29242
box 0 0 1 1
use contact_7  contact_7_107
timestamp 1624857261
transform 1 0 6041 0 1 29237
box 0 0 1 1
use and3_dec  and3_dec_53
timestamp 1624857261
transform 1 0 5803 0 1 29230
box 0 -60 2072 490
use contact_7  contact_7_432
timestamp 1624857261
transform 1 0 7676 0 1 26823
box 0 0 1 1
use contact_19  contact_19_432
timestamp 1624857261
transform 1 0 7677 0 1 26828
box 0 0 1 1
use contact_7  contact_7_435
timestamp 1624857261
transform 1 0 7676 0 1 26428
box 0 0 1 1
use contact_19  contact_19_435
timestamp 1624857261
transform 1 0 7677 0 1 26433
box 0 0 1 1
use contact_7  contact_7_426
timestamp 1624857261
transform 1 0 7676 0 1 27613
box 0 0 1 1
use contact_19  contact_19_426
timestamp 1624857261
transform 1 0 7677 0 1 27618
box 0 0 1 1
use contact_7  contact_7_429
timestamp 1624857261
transform 1 0 7676 0 1 27218
box 0 0 1 1
use contact_19  contact_19_429
timestamp 1624857261
transform 1 0 7677 0 1 27223
box 0 0 1 1
use contact_7  contact_7_417
timestamp 1624857261
transform 1 0 7676 0 1 28798
box 0 0 1 1
use contact_19  contact_19_417
timestamp 1624857261
transform 1 0 7677 0 1 28803
box 0 0 1 1
use contact_7  contact_7_420
timestamp 1624857261
transform 1 0 7676 0 1 28403
box 0 0 1 1
use contact_19  contact_19_420
timestamp 1624857261
transform 1 0 7677 0 1 28408
box 0 0 1 1
use contact_7  contact_7_423
timestamp 1624857261
transform 1 0 7676 0 1 28008
box 0 0 1 1
use contact_19  contact_19_423
timestamp 1624857261
transform 1 0 7677 0 1 28013
box 0 0 1 1
use contact_7  contact_7_414
timestamp 1624857261
transform 1 0 7676 0 1 29193
box 0 0 1 1
use contact_19  contact_19_414
timestamp 1624857261
transform 1 0 7677 0 1 29198
box 0 0 1 1
use contact_17  contact_17_156
timestamp 1624857261
transform 1 0 5464 0 1 29708
box 0 0 1 1
use contact_17  contact_17_159
timestamp 1624857261
transform 1 0 5464 0 1 29484
box 0 0 1 1
use contact_7  contact_7_105
timestamp 1624857261
transform 1 0 6041 0 1 29611
box 0 0 1 1
use contact_19  contact_19_105
timestamp 1624857261
transform 1 0 6042 0 1 29616
box 0 0 1 1
use contact_7  contact_7_412
timestamp 1624857261
transform 1 0 6466 0 1 29611
box 0 0 1 1
use contact_19  contact_19_412
timestamp 1624857261
transform 1 0 6467 0 1 29616
box 0 0 1 1
use contact_7  contact_7_410
timestamp 1624857261
transform 1 0 6898 0 1 29611
box 0 0 1 1
use contact_19  contact_19_410
timestamp 1624857261
transform 1 0 6899 0 1 29616
box 0 0 1 1
use contact_7  contact_7_104
timestamp 1624857261
transform 1 0 7280 0 1 29588
box 0 0 1 1
use contact_19  contact_19_104
timestamp 1624857261
transform 1 0 7281 0 1 29593
box 0 0 1 1
use contact_17  contact_17_158
timestamp 1624857261
transform 1 0 4744 0 1 29910
box 0 0 1 1
use contact_17  contact_17_157
timestamp 1624857261
transform 1 0 4984 0 1 29798
box 0 0 1 1
use contact_19  contact_19_409
timestamp 1624857261
transform 1 0 6467 0 1 29974
box 0 0 1 1
use contact_7  contact_7_409
timestamp 1624857261
transform 1 0 6466 0 1 29969
box 0 0 1 1
use contact_19  contact_19_407
timestamp 1624857261
transform 1 0 6899 0 1 29974
box 0 0 1 1
use contact_7  contact_7_407
timestamp 1624857261
transform 1 0 6898 0 1 29969
box 0 0 1 1
use contact_19  contact_19_102
timestamp 1624857261
transform 1 0 7281 0 1 29988
box 0 0 1 1
use contact_7  contact_7_102
timestamp 1624857261
transform 1 0 7280 0 1 29983
box 0 0 1 1
use and3_dec  and3_dec_52
timestamp 1624857261
transform 1 0 5803 0 -1 30020
box 0 -60 2072 490
use and3_dec  and3_dec_51
timestamp 1624857261
transform 1 0 5803 0 1 30020
box 0 -60 2072 490
use contact_17  contact_17_155
timestamp 1624857261
transform 1 0 4504 0 1 30072
box 0 0 1 1
use contact_17  contact_17_154
timestamp 1624857261
transform 1 0 5064 0 1 30184
box 0 0 1 1
use contact_17  contact_17_153
timestamp 1624857261
transform 1 0 5464 0 1 30274
box 0 0 1 1
use contact_19  contact_19_103
timestamp 1624857261
transform 1 0 6042 0 1 30032
box 0 0 1 1
use contact_7  contact_7_103
timestamp 1624857261
transform 1 0 6041 0 1 30027
box 0 0 1 1
use contact_17  contact_17_150
timestamp 1624857261
transform 1 0 5464 0 1 30498
box 0 0 1 1
use contact_19  contact_19_406
timestamp 1624857261
transform 1 0 6467 0 1 30406
box 0 0 1 1
use contact_7  contact_7_406
timestamp 1624857261
transform 1 0 6466 0 1 30401
box 0 0 1 1
use contact_19  contact_19_404
timestamp 1624857261
transform 1 0 6899 0 1 30406
box 0 0 1 1
use contact_7  contact_7_404
timestamp 1624857261
transform 1 0 6898 0 1 30401
box 0 0 1 1
use contact_19  contact_19_101
timestamp 1624857261
transform 1 0 6042 0 1 30406
box 0 0 1 1
use contact_7  contact_7_101
timestamp 1624857261
transform 1 0 6041 0 1 30401
box 0 0 1 1
use contact_19  contact_19_100
timestamp 1624857261
transform 1 0 7281 0 1 30383
box 0 0 1 1
use contact_7  contact_7_100
timestamp 1624857261
transform 1 0 7280 0 1 30378
box 0 0 1 1
use and3_dec  and3_dec_50
timestamp 1624857261
transform 1 0 5803 0 -1 30810
box 0 -60 2072 490
use contact_17  contact_17_152
timestamp 1624857261
transform 1 0 4584 0 1 30700
box 0 0 1 1
use contact_17  contact_17_151
timestamp 1624857261
transform 1 0 5064 0 1 30588
box 0 0 1 1
use contact_7  contact_7_99
timestamp 1624857261
transform 1 0 6041 0 1 30817
box 0 0 1 1
use contact_19  contact_19_99
timestamp 1624857261
transform 1 0 6042 0 1 30822
box 0 0 1 1
use contact_7  contact_7_403
timestamp 1624857261
transform 1 0 6466 0 1 30759
box 0 0 1 1
use contact_19  contact_19_403
timestamp 1624857261
transform 1 0 6467 0 1 30764
box 0 0 1 1
use contact_7  contact_7_401
timestamp 1624857261
transform 1 0 6898 0 1 30759
box 0 0 1 1
use contact_19  contact_19_401
timestamp 1624857261
transform 1 0 6899 0 1 30764
box 0 0 1 1
use contact_7  contact_7_98
timestamp 1624857261
transform 1 0 7280 0 1 30773
box 0 0 1 1
use contact_19  contact_19_98
timestamp 1624857261
transform 1 0 7281 0 1 30778
box 0 0 1 1
use contact_17  contact_17_149
timestamp 1624857261
transform 1 0 4664 0 1 30862
box 0 0 1 1
use contact_17  contact_17_148
timestamp 1624857261
transform 1 0 5064 0 1 30974
box 0 0 1 1
use contact_17  contact_17_147
timestamp 1624857261
transform 1 0 5464 0 1 31064
box 0 0 1 1
use and3_dec  and3_dec_49
timestamp 1624857261
transform 1 0 5803 0 1 30810
box 0 -60 2072 490
use and3_dec  and3_dec_48
timestamp 1624857261
transform 1 0 5803 0 -1 31600
box 0 -60 2072 490
use contact_17  contact_17_145
timestamp 1624857261
transform 1 0 5064 0 1 31378
box 0 0 1 1
use contact_17  contact_17_144
timestamp 1624857261
transform 1 0 5464 0 1 31288
box 0 0 1 1
use contact_7  contact_7_97
timestamp 1624857261
transform 1 0 6041 0 1 31191
box 0 0 1 1
use contact_19  contact_19_97
timestamp 1624857261
transform 1 0 6042 0 1 31196
box 0 0 1 1
use contact_7  contact_7_400
timestamp 1624857261
transform 1 0 6466 0 1 31191
box 0 0 1 1
use contact_19  contact_19_400
timestamp 1624857261
transform 1 0 6467 0 1 31196
box 0 0 1 1
use contact_7  contact_7_398
timestamp 1624857261
transform 1 0 6898 0 1 31191
box 0 0 1 1
use contact_19  contact_19_398
timestamp 1624857261
transform 1 0 6899 0 1 31196
box 0 0 1 1
use contact_7  contact_7_96
timestamp 1624857261
transform 1 0 7280 0 1 31168
box 0 0 1 1
use contact_19  contact_19_96
timestamp 1624857261
transform 1 0 7281 0 1 31173
box 0 0 1 1
use contact_17  contact_17_143
timestamp 1624857261
transform 1 0 4504 0 1 31652
box 0 0 1 1
use contact_17  contact_17_146
timestamp 1624857261
transform 1 0 4744 0 1 31490
box 0 0 1 1
use contact_7  contact_7_95
timestamp 1624857261
transform 1 0 6041 0 1 31607
box 0 0 1 1
use contact_19  contact_19_95
timestamp 1624857261
transform 1 0 6042 0 1 31612
box 0 0 1 1
use contact_7  contact_7_397
timestamp 1624857261
transform 1 0 6466 0 1 31549
box 0 0 1 1
use contact_19  contact_19_397
timestamp 1624857261
transform 1 0 6467 0 1 31554
box 0 0 1 1
use contact_7  contact_7_395
timestamp 1624857261
transform 1 0 6898 0 1 31549
box 0 0 1 1
use contact_19  contact_19_395
timestamp 1624857261
transform 1 0 6899 0 1 31554
box 0 0 1 1
use contact_7  contact_7_94
timestamp 1624857261
transform 1 0 7280 0 1 31563
box 0 0 1 1
use contact_19  contact_19_94
timestamp 1624857261
transform 1 0 7281 0 1 31568
box 0 0 1 1
use and3_dec  and3_dec_47
timestamp 1624857261
transform 1 0 5803 0 1 31600
box 0 -60 2072 490
use contact_17  contact_17_142
timestamp 1624857261
transform 1 0 4824 0 1 31764
box 0 0 1 1
use contact_17  contact_17_141
timestamp 1624857261
transform 1 0 5544 0 1 31854
box 0 0 1 1
use contact_17  contact_17_139
timestamp 1624857261
transform 1 0 4824 0 1 32168
box 0 0 1 1
use contact_17  contact_17_138
timestamp 1624857261
transform 1 0 5544 0 1 32078
box 0 0 1 1
use contact_7  contact_7_93
timestamp 1624857261
transform 1 0 6041 0 1 31981
box 0 0 1 1
use contact_19  contact_19_93
timestamp 1624857261
transform 1 0 6042 0 1 31986
box 0 0 1 1
use contact_7  contact_7_394
timestamp 1624857261
transform 1 0 6466 0 1 31981
box 0 0 1 1
use contact_19  contact_19_394
timestamp 1624857261
transform 1 0 6467 0 1 31986
box 0 0 1 1
use contact_7  contact_7_392
timestamp 1624857261
transform 1 0 6898 0 1 31981
box 0 0 1 1
use contact_19  contact_19_392
timestamp 1624857261
transform 1 0 6899 0 1 31986
box 0 0 1 1
use contact_7  contact_7_92
timestamp 1624857261
transform 1 0 7280 0 1 31958
box 0 0 1 1
use contact_19  contact_19_92
timestamp 1624857261
transform 1 0 7281 0 1 31963
box 0 0 1 1
use and3_dec  and3_dec_46
timestamp 1624857261
transform 1 0 5803 0 -1 32390
box 0 -60 2072 490
use contact_17  contact_17_137
timestamp 1624857261
transform 1 0 4664 0 1 32442
box 0 0 1 1
use contact_17  contact_17_140
timestamp 1624857261
transform 1 0 4584 0 1 32280
box 0 0 1 1
use contact_7  contact_7_91
timestamp 1624857261
transform 1 0 6041 0 1 32397
box 0 0 1 1
use contact_19  contact_19_91
timestamp 1624857261
transform 1 0 6042 0 1 32402
box 0 0 1 1
use contact_7  contact_7_391
timestamp 1624857261
transform 1 0 6466 0 1 32339
box 0 0 1 1
use contact_19  contact_19_391
timestamp 1624857261
transform 1 0 6467 0 1 32344
box 0 0 1 1
use contact_7  contact_7_389
timestamp 1624857261
transform 1 0 6898 0 1 32339
box 0 0 1 1
use contact_19  contact_19_389
timestamp 1624857261
transform 1 0 6899 0 1 32344
box 0 0 1 1
use contact_7  contact_7_90
timestamp 1624857261
transform 1 0 7280 0 1 32353
box 0 0 1 1
use contact_19  contact_19_90
timestamp 1624857261
transform 1 0 7281 0 1 32358
box 0 0 1 1
use contact_17  contact_17_136
timestamp 1624857261
transform 1 0 4824 0 1 32554
box 0 0 1 1
use contact_17  contact_17_135
timestamp 1624857261
transform 1 0 5544 0 1 32644
box 0 0 1 1
use contact_7  contact_7_88
timestamp 1624857261
transform 1 0 7280 0 1 32748
box 0 0 1 1
use and3_dec  and3_dec_45
timestamp 1624857261
transform 1 0 5803 0 1 32390
box 0 -60 2072 490
use and3_dec  and3_dec_44
timestamp 1624857261
transform 1 0 5803 0 -1 33180
box 0 -60 2072 490
use contact_7  contact_7_408
timestamp 1624857261
transform 1 0 7676 0 1 29983
box 0 0 1 1
use contact_19  contact_19_408
timestamp 1624857261
transform 1 0 7677 0 1 29988
box 0 0 1 1
use contact_7  contact_7_411
timestamp 1624857261
transform 1 0 7676 0 1 29588
box 0 0 1 1
use contact_19  contact_19_411
timestamp 1624857261
transform 1 0 7677 0 1 29593
box 0 0 1 1
use contact_7  contact_7_399
timestamp 1624857261
transform 1 0 7676 0 1 31168
box 0 0 1 1
use contact_19  contact_19_399
timestamp 1624857261
transform 1 0 7677 0 1 31173
box 0 0 1 1
use contact_7  contact_7_402
timestamp 1624857261
transform 1 0 7676 0 1 30773
box 0 0 1 1
use contact_19  contact_19_402
timestamp 1624857261
transform 1 0 7677 0 1 30778
box 0 0 1 1
use contact_7  contact_7_405
timestamp 1624857261
transform 1 0 7676 0 1 30378
box 0 0 1 1
use contact_19  contact_19_405
timestamp 1624857261
transform 1 0 7677 0 1 30383
box 0 0 1 1
use contact_7  contact_7_393
timestamp 1624857261
transform 1 0 7676 0 1 31958
box 0 0 1 1
use contact_19  contact_19_393
timestamp 1624857261
transform 1 0 7677 0 1 31963
box 0 0 1 1
use contact_7  contact_7_396
timestamp 1624857261
transform 1 0 7676 0 1 31563
box 0 0 1 1
use contact_19  contact_19_396
timestamp 1624857261
transform 1 0 7677 0 1 31568
box 0 0 1 1
use contact_7  contact_7_387
timestamp 1624857261
transform 1 0 7676 0 1 32748
box 0 0 1 1
use contact_7  contact_7_390
timestamp 1624857261
transform 1 0 7676 0 1 32353
box 0 0 1 1
use contact_19  contact_19_390
timestamp 1624857261
transform 1 0 7677 0 1 32358
box 0 0 1 1
use contact_17  contact_17_133
timestamp 1624857261
transform 1 0 4824 0 1 32958
box 0 0 1 1
use contact_17  contact_17_132
timestamp 1624857261
transform 1 0 5544 0 1 32868
box 0 0 1 1
use contact_19  contact_19_388
timestamp 1624857261
transform 1 0 6467 0 1 32776
box 0 0 1 1
use contact_7  contact_7_388
timestamp 1624857261
transform 1 0 6466 0 1 32771
box 0 0 1 1
use contact_19  contact_19_386
timestamp 1624857261
transform 1 0 6899 0 1 32776
box 0 0 1 1
use contact_7  contact_7_386
timestamp 1624857261
transform 1 0 6898 0 1 32771
box 0 0 1 1
use contact_19  contact_19_89
timestamp 1624857261
transform 1 0 6042 0 1 32776
box 0 0 1 1
use contact_7  contact_7_89
timestamp 1624857261
transform 1 0 6041 0 1 32771
box 0 0 1 1
use contact_19  contact_19_88
timestamp 1624857261
transform 1 0 7281 0 1 32753
box 0 0 1 1
use contact_17  contact_17_131
timestamp 1624857261
transform 1 0 4504 0 1 33232
box 0 0 1 1
use contact_17  contact_17_134
timestamp 1624857261
transform 1 0 4744 0 1 33070
box 0 0 1 1
use contact_7  contact_7_87
timestamp 1624857261
transform 1 0 6041 0 1 33187
box 0 0 1 1
use contact_19  contact_19_87
timestamp 1624857261
transform 1 0 6042 0 1 33192
box 0 0 1 1
use contact_7  contact_7_385
timestamp 1624857261
transform 1 0 6466 0 1 33129
box 0 0 1 1
use contact_19  contact_19_385
timestamp 1624857261
transform 1 0 6467 0 1 33134
box 0 0 1 1
use contact_7  contact_7_383
timestamp 1624857261
transform 1 0 6898 0 1 33129
box 0 0 1 1
use contact_19  contact_19_383
timestamp 1624857261
transform 1 0 6899 0 1 33134
box 0 0 1 1
use contact_7  contact_7_86
timestamp 1624857261
transform 1 0 7280 0 1 33143
box 0 0 1 1
use contact_19  contact_19_86
timestamp 1624857261
transform 1 0 7281 0 1 33148
box 0 0 1 1
use and3_dec  and3_dec_43
timestamp 1624857261
transform 1 0 5803 0 1 33180
box 0 -60 2072 490
use contact_17  contact_17_130
timestamp 1624857261
transform 1 0 4904 0 1 33344
box 0 0 1 1
use contact_17  contact_17_129
timestamp 1624857261
transform 1 0 5544 0 1 33434
box 0 0 1 1
use contact_7  contact_7_85
timestamp 1624857261
transform 1 0 6041 0 1 33561
box 0 0 1 1
use contact_19  contact_19_85
timestamp 1624857261
transform 1 0 6042 0 1 33566
box 0 0 1 1
use contact_7  contact_7_382
timestamp 1624857261
transform 1 0 6466 0 1 33561
box 0 0 1 1
use contact_19  contact_19_382
timestamp 1624857261
transform 1 0 6467 0 1 33566
box 0 0 1 1
use contact_7  contact_7_380
timestamp 1624857261
transform 1 0 6898 0 1 33561
box 0 0 1 1
use contact_19  contact_19_380
timestamp 1624857261
transform 1 0 6899 0 1 33566
box 0 0 1 1
use contact_7  contact_7_84
timestamp 1624857261
transform 1 0 7280 0 1 33538
box 0 0 1 1
use contact_19  contact_19_84
timestamp 1624857261
transform 1 0 7281 0 1 33543
box 0 0 1 1
use contact_17  contact_17_127
timestamp 1624857261
transform 1 0 4904 0 1 33748
box 0 0 1 1
use contact_17  contact_17_126
timestamp 1624857261
transform 1 0 5544 0 1 33658
box 0 0 1 1
use and3_dec  and3_dec_42
timestamp 1624857261
transform 1 0 5803 0 -1 33970
box 0 -60 2072 490
use contact_17  contact_17_125
timestamp 1624857261
transform 1 0 4664 0 1 34022
box 0 0 1 1
use contact_17  contact_17_128
timestamp 1624857261
transform 1 0 4584 0 1 33860
box 0 0 1 1
use contact_7  contact_7_83
timestamp 1624857261
transform 1 0 6041 0 1 33977
box 0 0 1 1
use contact_19  contact_19_83
timestamp 1624857261
transform 1 0 6042 0 1 33982
box 0 0 1 1
use contact_7  contact_7_379
timestamp 1624857261
transform 1 0 6466 0 1 33919
box 0 0 1 1
use contact_19  contact_19_379
timestamp 1624857261
transform 1 0 6467 0 1 33924
box 0 0 1 1
use contact_7  contact_7_377
timestamp 1624857261
transform 1 0 6898 0 1 33919
box 0 0 1 1
use contact_19  contact_19_377
timestamp 1624857261
transform 1 0 6899 0 1 33924
box 0 0 1 1
use contact_7  contact_7_82
timestamp 1624857261
transform 1 0 7280 0 1 33933
box 0 0 1 1
use contact_19  contact_19_82
timestamp 1624857261
transform 1 0 7281 0 1 33938
box 0 0 1 1
use contact_17  contact_17_124
timestamp 1624857261
transform 1 0 4904 0 1 34134
box 0 0 1 1
use contact_17  contact_17_123
timestamp 1624857261
transform 1 0 5544 0 1 34224
box 0 0 1 1
use contact_7  contact_7_81
timestamp 1624857261
transform 1 0 6041 0 1 34351
box 0 0 1 1
use contact_19  contact_19_81
timestamp 1624857261
transform 1 0 6042 0 1 34356
box 0 0 1 1
use contact_7  contact_7_376
timestamp 1624857261
transform 1 0 6466 0 1 34351
box 0 0 1 1
use contact_19  contact_19_376
timestamp 1624857261
transform 1 0 6467 0 1 34356
box 0 0 1 1
use contact_7  contact_7_374
timestamp 1624857261
transform 1 0 6898 0 1 34351
box 0 0 1 1
use contact_19  contact_19_374
timestamp 1624857261
transform 1 0 6899 0 1 34356
box 0 0 1 1
use contact_7  contact_7_80
timestamp 1624857261
transform 1 0 7280 0 1 34328
box 0 0 1 1
use contact_19  contact_19_80
timestamp 1624857261
transform 1 0 7281 0 1 34333
box 0 0 1 1
use and3_dec  and3_dec_41
timestamp 1624857261
transform 1 0 5803 0 1 33970
box 0 -60 2072 490
use and3_dec  and3_dec_40
timestamp 1624857261
transform 1 0 5803 0 -1 34760
box 0 -60 2072 490
use contact_17  contact_17_122
timestamp 1624857261
transform 1 0 4744 0 1 34650
box 0 0 1 1
use contact_17  contact_17_121
timestamp 1624857261
transform 1 0 4904 0 1 34538
box 0 0 1 1
use contact_17  contact_17_120
timestamp 1624857261
transform 1 0 5544 0 1 34448
box 0 0 1 1
use contact_17  contact_17_119
timestamp 1624857261
transform 1 0 4504 0 1 34812
box 0 0 1 1
use contact_17  contact_17_118
timestamp 1624857261
transform 1 0 4984 0 1 34924
box 0 0 1 1
use contact_7  contact_7_79
timestamp 1624857261
transform 1 0 6041 0 1 34767
box 0 0 1 1
use contact_19  contact_19_79
timestamp 1624857261
transform 1 0 6042 0 1 34772
box 0 0 1 1
use contact_7  contact_7_373
timestamp 1624857261
transform 1 0 6466 0 1 34709
box 0 0 1 1
use contact_19  contact_19_373
timestamp 1624857261
transform 1 0 6467 0 1 34714
box 0 0 1 1
use contact_7  contact_7_371
timestamp 1624857261
transform 1 0 6898 0 1 34709
box 0 0 1 1
use contact_19  contact_19_371
timestamp 1624857261
transform 1 0 6899 0 1 34714
box 0 0 1 1
use contact_7  contact_7_78
timestamp 1624857261
transform 1 0 7280 0 1 34723
box 0 0 1 1
use contact_19  contact_19_78
timestamp 1624857261
transform 1 0 7281 0 1 34728
box 0 0 1 1
use and3_dec  and3_dec_39
timestamp 1624857261
transform 1 0 5803 0 1 34760
box 0 -60 2072 490
use contact_17  contact_17_117
timestamp 1624857261
transform 1 0 5544 0 1 35014
box 0 0 1 1
use contact_19  contact_19_370
timestamp 1624857261
transform 1 0 6467 0 1 35146
box 0 0 1 1
use contact_7  contact_7_370
timestamp 1624857261
transform 1 0 6466 0 1 35141
box 0 0 1 1
use contact_19  contact_19_368
timestamp 1624857261
transform 1 0 6899 0 1 35146
box 0 0 1 1
use contact_7  contact_7_368
timestamp 1624857261
transform 1 0 6898 0 1 35141
box 0 0 1 1
use contact_19  contact_19_77
timestamp 1624857261
transform 1 0 6042 0 1 35146
box 0 0 1 1
use contact_7  contact_7_77
timestamp 1624857261
transform 1 0 6041 0 1 35141
box 0 0 1 1
use contact_19  contact_19_76
timestamp 1624857261
transform 1 0 7281 0 1 35123
box 0 0 1 1
use contact_7  contact_7_76
timestamp 1624857261
transform 1 0 7280 0 1 35118
box 0 0 1 1
use contact_17  contact_17_116
timestamp 1624857261
transform 1 0 4584 0 1 35440
box 0 0 1 1
use contact_17  contact_17_115
timestamp 1624857261
transform 1 0 4984 0 1 35328
box 0 0 1 1
use contact_17  contact_17_114
timestamp 1624857261
transform 1 0 5544 0 1 35238
box 0 0 1 1
use contact_19  contact_19_367
timestamp 1624857261
transform 1 0 6467 0 1 35504
box 0 0 1 1
use contact_7  contact_7_367
timestamp 1624857261
transform 1 0 6466 0 1 35499
box 0 0 1 1
use contact_19  contact_19_365
timestamp 1624857261
transform 1 0 6899 0 1 35504
box 0 0 1 1
use contact_7  contact_7_365
timestamp 1624857261
transform 1 0 6898 0 1 35499
box 0 0 1 1
use and3_dec  and3_dec_38
timestamp 1624857261
transform 1 0 5803 0 -1 35550
box 0 -60 2072 490
use and3_dec  and3_dec_37
timestamp 1624857261
transform 1 0 5803 0 1 35550
box 0 -60 2072 490
use contact_17  contact_17_113
timestamp 1624857261
transform 1 0 4664 0 1 35602
box 0 0 1 1
use contact_17  contact_17_112
timestamp 1624857261
transform 1 0 4984 0 1 35714
box 0 0 1 1
use contact_19  contact_19_75
timestamp 1624857261
transform 1 0 6042 0 1 35562
box 0 0 1 1
use contact_7  contact_7_75
timestamp 1624857261
transform 1 0 6041 0 1 35557
box 0 0 1 1
use contact_19  contact_19_74
timestamp 1624857261
transform 1 0 7281 0 1 35518
box 0 0 1 1
use contact_7  contact_7_74
timestamp 1624857261
transform 1 0 7280 0 1 35513
box 0 0 1 1
use contact_17  contact_17_108
timestamp 1624857261
transform 1 0 5544 0 1 36028
box 0 0 1 1
use contact_17  contact_17_111
timestamp 1624857261
transform 1 0 5544 0 1 35804
box 0 0 1 1
use contact_7  contact_7_73
timestamp 1624857261
transform 1 0 6041 0 1 35931
box 0 0 1 1
use contact_19  contact_19_73
timestamp 1624857261
transform 1 0 6042 0 1 35936
box 0 0 1 1
use contact_7  contact_7_364
timestamp 1624857261
transform 1 0 6466 0 1 35931
box 0 0 1 1
use contact_19  contact_19_364
timestamp 1624857261
transform 1 0 6467 0 1 35936
box 0 0 1 1
use contact_7  contact_7_362
timestamp 1624857261
transform 1 0 6898 0 1 35931
box 0 0 1 1
use contact_19  contact_19_362
timestamp 1624857261
transform 1 0 6899 0 1 35936
box 0 0 1 1
use contact_7  contact_7_72
timestamp 1624857261
transform 1 0 7280 0 1 35908
box 0 0 1 1
use contact_19  contact_19_72
timestamp 1624857261
transform 1 0 7281 0 1 35913
box 0 0 1 1
use and3_dec  and3_dec_36
timestamp 1624857261
transform 1 0 5803 0 -1 36340
box 0 -60 2072 490
use contact_7  contact_7_381
timestamp 1624857261
transform 1 0 7676 0 1 33538
box 0 0 1 1
use contact_19  contact_19_381
timestamp 1624857261
transform 1 0 7677 0 1 33543
box 0 0 1 1
use contact_7  contact_7_384
timestamp 1624857261
transform 1 0 7676 0 1 33143
box 0 0 1 1
use contact_19  contact_19_384
timestamp 1624857261
transform 1 0 7677 0 1 33148
box 0 0 1 1
use contact_19  contact_19_387
timestamp 1624857261
transform 1 0 7677 0 1 32753
box 0 0 1 1
use contact_7  contact_7_375
timestamp 1624857261
transform 1 0 7676 0 1 34328
box 0 0 1 1
use contact_19  contact_19_375
timestamp 1624857261
transform 1 0 7677 0 1 34333
box 0 0 1 1
use contact_7  contact_7_378
timestamp 1624857261
transform 1 0 7676 0 1 33933
box 0 0 1 1
use contact_19  contact_19_378
timestamp 1624857261
transform 1 0 7677 0 1 33938
box 0 0 1 1
use contact_7  contact_7_369
timestamp 1624857261
transform 1 0 7676 0 1 35118
box 0 0 1 1
use contact_19  contact_19_369
timestamp 1624857261
transform 1 0 7677 0 1 35123
box 0 0 1 1
use contact_7  contact_7_372
timestamp 1624857261
transform 1 0 7676 0 1 34723
box 0 0 1 1
use contact_19  contact_19_372
timestamp 1624857261
transform 1 0 7677 0 1 34728
box 0 0 1 1
use contact_7  contact_7_363
timestamp 1624857261
transform 1 0 7676 0 1 35908
box 0 0 1 1
use contact_19  contact_19_363
timestamp 1624857261
transform 1 0 7677 0 1 35913
box 0 0 1 1
use contact_7  contact_7_366
timestamp 1624857261
transform 1 0 7676 0 1 35513
box 0 0 1 1
use contact_19  contact_19_366
timestamp 1624857261
transform 1 0 7677 0 1 35518
box 0 0 1 1
use contact_17  contact_17_110
timestamp 1624857261
transform 1 0 4744 0 1 36230
box 0 0 1 1
use contact_17  contact_17_109
timestamp 1624857261
transform 1 0 4984 0 1 36118
box 0 0 1 1
use contact_19  contact_19_361
timestamp 1624857261
transform 1 0 6467 0 1 36294
box 0 0 1 1
use contact_7  contact_7_361
timestamp 1624857261
transform 1 0 6466 0 1 36289
box 0 0 1 1
use contact_19  contact_19_359
timestamp 1624857261
transform 1 0 6899 0 1 36294
box 0 0 1 1
use contact_7  contact_7_359
timestamp 1624857261
transform 1 0 6898 0 1 36289
box 0 0 1 1
use contact_7  contact_7_70
timestamp 1624857261
transform 1 0 7280 0 1 36303
box 0 0 1 1
use contact_17  contact_17_107
timestamp 1624857261
transform 1 0 4504 0 1 36392
box 0 0 1 1
use contact_17  contact_17_106
timestamp 1624857261
transform 1 0 5064 0 1 36504
box 0 0 1 1
use contact_19  contact_19_71
timestamp 1624857261
transform 1 0 6042 0 1 36352
box 0 0 1 1
use contact_7  contact_7_71
timestamp 1624857261
transform 1 0 6041 0 1 36347
box 0 0 1 1
use contact_19  contact_19_70
timestamp 1624857261
transform 1 0 7281 0 1 36308
box 0 0 1 1
use and3_dec  and3_dec_35
timestamp 1624857261
transform 1 0 5803 0 1 36340
box 0 -60 2072 490
use contact_17  contact_17_102
timestamp 1624857261
transform 1 0 5544 0 1 36818
box 0 0 1 1
use contact_17  contact_17_105
timestamp 1624857261
transform 1 0 5544 0 1 36594
box 0 0 1 1
use contact_7  contact_7_69
timestamp 1624857261
transform 1 0 6041 0 1 36721
box 0 0 1 1
use contact_19  contact_19_69
timestamp 1624857261
transform 1 0 6042 0 1 36726
box 0 0 1 1
use contact_7  contact_7_358
timestamp 1624857261
transform 1 0 6466 0 1 36721
box 0 0 1 1
use contact_19  contact_19_358
timestamp 1624857261
transform 1 0 6467 0 1 36726
box 0 0 1 1
use contact_7  contact_7_356
timestamp 1624857261
transform 1 0 6898 0 1 36721
box 0 0 1 1
use contact_19  contact_19_356
timestamp 1624857261
transform 1 0 6899 0 1 36726
box 0 0 1 1
use contact_7  contact_7_68
timestamp 1624857261
transform 1 0 7280 0 1 36698
box 0 0 1 1
use contact_19  contact_19_68
timestamp 1624857261
transform 1 0 7281 0 1 36703
box 0 0 1 1
use contact_17  contact_17_104
timestamp 1624857261
transform 1 0 4584 0 1 37020
box 0 0 1 1
use contact_17  contact_17_103
timestamp 1624857261
transform 1 0 5064 0 1 36908
box 0 0 1 1
use contact_19  contact_19_355
timestamp 1624857261
transform 1 0 6467 0 1 37084
box 0 0 1 1
use contact_7  contact_7_355
timestamp 1624857261
transform 1 0 6466 0 1 37079
box 0 0 1 1
use contact_19  contact_19_353
timestamp 1624857261
transform 1 0 6899 0 1 37084
box 0 0 1 1
use contact_7  contact_7_353
timestamp 1624857261
transform 1 0 6898 0 1 37079
box 0 0 1 1
use contact_19  contact_19_66
timestamp 1624857261
transform 1 0 7281 0 1 37098
box 0 0 1 1
use contact_7  contact_7_66
timestamp 1624857261
transform 1 0 7280 0 1 37093
box 0 0 1 1
use and3_dec  and3_dec_34
timestamp 1624857261
transform 1 0 5803 0 -1 37130
box 0 -60 2072 490
use and3_dec  and3_dec_33
timestamp 1624857261
transform 1 0 5803 0 1 37130
box 0 -60 2072 490
use contact_17  contact_17_101
timestamp 1624857261
transform 1 0 4664 0 1 37182
box 0 0 1 1
use contact_17  contact_17_100
timestamp 1624857261
transform 1 0 5064 0 1 37294
box 0 0 1 1
use contact_17  contact_17_99
timestamp 1624857261
transform 1 0 5544 0 1 37384
box 0 0 1 1
use contact_19  contact_19_67
timestamp 1624857261
transform 1 0 6042 0 1 37142
box 0 0 1 1
use contact_7  contact_7_67
timestamp 1624857261
transform 1 0 6041 0 1 37137
box 0 0 1 1
use contact_17  contact_17_96
timestamp 1624857261
transform 1 0 5544 0 1 37608
box 0 0 1 1
use contact_19  contact_19_352
timestamp 1624857261
transform 1 0 6467 0 1 37516
box 0 0 1 1
use contact_7  contact_7_352
timestamp 1624857261
transform 1 0 6466 0 1 37511
box 0 0 1 1
use contact_19  contact_19_350
timestamp 1624857261
transform 1 0 6899 0 1 37516
box 0 0 1 1
use contact_7  contact_7_350
timestamp 1624857261
transform 1 0 6898 0 1 37511
box 0 0 1 1
use contact_19  contact_19_65
timestamp 1624857261
transform 1 0 6042 0 1 37516
box 0 0 1 1
use contact_7  contact_7_65
timestamp 1624857261
transform 1 0 6041 0 1 37511
box 0 0 1 1
use contact_19  contact_19_64
timestamp 1624857261
transform 1 0 7281 0 1 37493
box 0 0 1 1
use contact_7  contact_7_64
timestamp 1624857261
transform 1 0 7280 0 1 37488
box 0 0 1 1
use and3_dec  and3_dec_32
timestamp 1624857261
transform 1 0 5803 0 -1 37920
box 0 -60 2072 490
use contact_17  contact_17_98
timestamp 1624857261
transform 1 0 4744 0 1 37810
box 0 0 1 1
use contact_17  contact_17_97
timestamp 1624857261
transform 1 0 5064 0 1 37698
box 0 0 1 1
use contact_7  contact_7_63
timestamp 1624857261
transform 1 0 6041 0 1 37927
box 0 0 1 1
use contact_19  contact_19_63
timestamp 1624857261
transform 1 0 6042 0 1 37932
box 0 0 1 1
use contact_7  contact_7_349
timestamp 1624857261
transform 1 0 6466 0 1 37869
box 0 0 1 1
use contact_19  contact_19_349
timestamp 1624857261
transform 1 0 6467 0 1 37874
box 0 0 1 1
use contact_7  contact_7_347
timestamp 1624857261
transform 1 0 6898 0 1 37869
box 0 0 1 1
use contact_19  contact_19_347
timestamp 1624857261
transform 1 0 6899 0 1 37874
box 0 0 1 1
use contact_7  contact_7_62
timestamp 1624857261
transform 1 0 7280 0 1 37883
box 0 0 1 1
use contact_19  contact_19_62
timestamp 1624857261
transform 1 0 7281 0 1 37888
box 0 0 1 1
use contact_17  contact_17_95
timestamp 1624857261
transform 1 0 4504 0 1 37972
box 0 0 1 1
use contact_17  contact_17_94
timestamp 1624857261
transform 1 0 4824 0 1 38084
box 0 0 1 1
use contact_17  contact_17_93
timestamp 1624857261
transform 1 0 5624 0 1 38174
box 0 0 1 1
use and3_dec  and3_dec_31
timestamp 1624857261
transform 1 0 5803 0 1 37920
box 0 -60 2072 490
use and3_dec  and3_dec_30
timestamp 1624857261
transform 1 0 5803 0 -1 38710
box 0 -60 2072 490
use contact_17  contact_17_91
timestamp 1624857261
transform 1 0 4824 0 1 38488
box 0 0 1 1
use contact_17  contact_17_90
timestamp 1624857261
transform 1 0 5624 0 1 38398
box 0 0 1 1
use contact_7  contact_7_61
timestamp 1624857261
transform 1 0 6041 0 1 38301
box 0 0 1 1
use contact_19  contact_19_61
timestamp 1624857261
transform 1 0 6042 0 1 38306
box 0 0 1 1
use contact_7  contact_7_346
timestamp 1624857261
transform 1 0 6466 0 1 38301
box 0 0 1 1
use contact_19  contact_19_346
timestamp 1624857261
transform 1 0 6467 0 1 38306
box 0 0 1 1
use contact_7  contact_7_344
timestamp 1624857261
transform 1 0 6898 0 1 38301
box 0 0 1 1
use contact_19  contact_19_344
timestamp 1624857261
transform 1 0 6899 0 1 38306
box 0 0 1 1
use contact_7  contact_7_60
timestamp 1624857261
transform 1 0 7280 0 1 38278
box 0 0 1 1
use contact_19  contact_19_60
timestamp 1624857261
transform 1 0 7281 0 1 38283
box 0 0 1 1
use contact_17  contact_17_89
timestamp 1624857261
transform 1 0 4664 0 1 38762
box 0 0 1 1
use contact_17  contact_17_92
timestamp 1624857261
transform 1 0 4584 0 1 38600
box 0 0 1 1
use contact_7  contact_7_59
timestamp 1624857261
transform 1 0 6041 0 1 38717
box 0 0 1 1
use contact_19  contact_19_59
timestamp 1624857261
transform 1 0 6042 0 1 38722
box 0 0 1 1
use contact_7  contact_7_343
timestamp 1624857261
transform 1 0 6466 0 1 38659
box 0 0 1 1
use contact_19  contact_19_343
timestamp 1624857261
transform 1 0 6467 0 1 38664
box 0 0 1 1
use contact_7  contact_7_341
timestamp 1624857261
transform 1 0 6898 0 1 38659
box 0 0 1 1
use contact_19  contact_19_341
timestamp 1624857261
transform 1 0 6899 0 1 38664
box 0 0 1 1
use contact_7  contact_7_58
timestamp 1624857261
transform 1 0 7280 0 1 38673
box 0 0 1 1
use contact_19  contact_19_58
timestamp 1624857261
transform 1 0 7281 0 1 38678
box 0 0 1 1
use and3_dec  and3_dec_29
timestamp 1624857261
transform 1 0 5803 0 1 38710
box 0 -60 2072 490
use contact_17  contact_17_88
timestamp 1624857261
transform 1 0 4824 0 1 38874
box 0 0 1 1
use contact_17  contact_17_87
timestamp 1624857261
transform 1 0 5624 0 1 38964
box 0 0 1 1
use contact_17  contact_17_85
timestamp 1624857261
transform 1 0 4824 0 1 39278
box 0 0 1 1
use contact_17  contact_17_84
timestamp 1624857261
transform 1 0 5624 0 1 39188
box 0 0 1 1
use contact_7  contact_7_57
timestamp 1624857261
transform 1 0 6041 0 1 39091
box 0 0 1 1
use contact_19  contact_19_57
timestamp 1624857261
transform 1 0 6042 0 1 39096
box 0 0 1 1
use contact_7  contact_7_340
timestamp 1624857261
transform 1 0 6466 0 1 39091
box 0 0 1 1
use contact_19  contact_19_340
timestamp 1624857261
transform 1 0 6467 0 1 39096
box 0 0 1 1
use contact_7  contact_7_338
timestamp 1624857261
transform 1 0 6898 0 1 39091
box 0 0 1 1
use contact_19  contact_19_338
timestamp 1624857261
transform 1 0 6899 0 1 39096
box 0 0 1 1
use contact_7  contact_7_56
timestamp 1624857261
transform 1 0 7280 0 1 39068
box 0 0 1 1
use contact_19  contact_19_56
timestamp 1624857261
transform 1 0 7281 0 1 39073
box 0 0 1 1
use and3_dec  and3_dec_28
timestamp 1624857261
transform 1 0 5803 0 -1 39500
box 0 -60 2072 490
use contact_7  contact_7_357
timestamp 1624857261
transform 1 0 7676 0 1 36698
box 0 0 1 1
use contact_19  contact_19_357
timestamp 1624857261
transform 1 0 7677 0 1 36703
box 0 0 1 1
use contact_7  contact_7_360
timestamp 1624857261
transform 1 0 7676 0 1 36303
box 0 0 1 1
use contact_19  contact_19_360
timestamp 1624857261
transform 1 0 7677 0 1 36308
box 0 0 1 1
use contact_7  contact_7_351
timestamp 1624857261
transform 1 0 7676 0 1 37488
box 0 0 1 1
use contact_19  contact_19_351
timestamp 1624857261
transform 1 0 7677 0 1 37493
box 0 0 1 1
use contact_7  contact_7_354
timestamp 1624857261
transform 1 0 7676 0 1 37093
box 0 0 1 1
use contact_19  contact_19_354
timestamp 1624857261
transform 1 0 7677 0 1 37098
box 0 0 1 1
use contact_7  contact_7_342
timestamp 1624857261
transform 1 0 7676 0 1 38673
box 0 0 1 1
use contact_7  contact_7_345
timestamp 1624857261
transform 1 0 7676 0 1 38278
box 0 0 1 1
use contact_19  contact_19_345
timestamp 1624857261
transform 1 0 7677 0 1 38283
box 0 0 1 1
use contact_7  contact_7_348
timestamp 1624857261
transform 1 0 7676 0 1 37883
box 0 0 1 1
use contact_19  contact_19_348
timestamp 1624857261
transform 1 0 7677 0 1 37888
box 0 0 1 1
use contact_7  contact_7_339
timestamp 1624857261
transform 1 0 7676 0 1 39068
box 0 0 1 1
use contact_19  contact_19_339
timestamp 1624857261
transform 1 0 7677 0 1 39073
box 0 0 1 1
use contact_19  contact_19_342
timestamp 1624857261
transform 1 0 7677 0 1 38678
box 0 0 1 1
use contact_17  contact_17_83
timestamp 1624857261
transform 1 0 4504 0 1 39552
box 0 0 1 1
use contact_17  contact_17_86
timestamp 1624857261
transform 1 0 4744 0 1 39390
box 0 0 1 1
use contact_7  contact_7_55
timestamp 1624857261
transform 1 0 6041 0 1 39507
box 0 0 1 1
use contact_19  contact_19_55
timestamp 1624857261
transform 1 0 6042 0 1 39512
box 0 0 1 1
use contact_7  contact_7_337
timestamp 1624857261
transform 1 0 6466 0 1 39449
box 0 0 1 1
use contact_19  contact_19_337
timestamp 1624857261
transform 1 0 6467 0 1 39454
box 0 0 1 1
use contact_7  contact_7_335
timestamp 1624857261
transform 1 0 6898 0 1 39449
box 0 0 1 1
use contact_19  contact_19_335
timestamp 1624857261
transform 1 0 6899 0 1 39454
box 0 0 1 1
use contact_7  contact_7_54
timestamp 1624857261
transform 1 0 7280 0 1 39463
box 0 0 1 1
use contact_19  contact_19_54
timestamp 1624857261
transform 1 0 7281 0 1 39468
box 0 0 1 1
use contact_17  contact_17_82
timestamp 1624857261
transform 1 0 4904 0 1 39664
box 0 0 1 1
use contact_17  contact_17_81
timestamp 1624857261
transform 1 0 5624 0 1 39754
box 0 0 1 1
use contact_7  contact_7_52
timestamp 1624857261
transform 1 0 7280 0 1 39858
box 0 0 1 1
use and3_dec  and3_dec_27
timestamp 1624857261
transform 1 0 5803 0 1 39500
box 0 -60 2072 490
use and3_dec  and3_dec_26
timestamp 1624857261
transform 1 0 5803 0 -1 40290
box 0 -60 2072 490
use contact_17  contact_17_79
timestamp 1624857261
transform 1 0 4904 0 1 40068
box 0 0 1 1
use contact_17  contact_17_78
timestamp 1624857261
transform 1 0 5624 0 1 39978
box 0 0 1 1
use contact_19  contact_19_334
timestamp 1624857261
transform 1 0 6467 0 1 39886
box 0 0 1 1
use contact_7  contact_7_334
timestamp 1624857261
transform 1 0 6466 0 1 39881
box 0 0 1 1
use contact_19  contact_19_332
timestamp 1624857261
transform 1 0 6899 0 1 39886
box 0 0 1 1
use contact_7  contact_7_332
timestamp 1624857261
transform 1 0 6898 0 1 39881
box 0 0 1 1
use contact_19  contact_19_53
timestamp 1624857261
transform 1 0 6042 0 1 39886
box 0 0 1 1
use contact_7  contact_7_53
timestamp 1624857261
transform 1 0 6041 0 1 39881
box 0 0 1 1
use contact_19  contact_19_52
timestamp 1624857261
transform 1 0 7281 0 1 39863
box 0 0 1 1
use contact_17  contact_17_77
timestamp 1624857261
transform 1 0 4664 0 1 40342
box 0 0 1 1
use contact_17  contact_17_80
timestamp 1624857261
transform 1 0 4584 0 1 40180
box 0 0 1 1
use contact_7  contact_7_51
timestamp 1624857261
transform 1 0 6041 0 1 40297
box 0 0 1 1
use contact_19  contact_19_51
timestamp 1624857261
transform 1 0 6042 0 1 40302
box 0 0 1 1
use contact_7  contact_7_331
timestamp 1624857261
transform 1 0 6466 0 1 40239
box 0 0 1 1
use contact_19  contact_19_331
timestamp 1624857261
transform 1 0 6467 0 1 40244
box 0 0 1 1
use contact_7  contact_7_329
timestamp 1624857261
transform 1 0 6898 0 1 40239
box 0 0 1 1
use contact_19  contact_19_329
timestamp 1624857261
transform 1 0 6899 0 1 40244
box 0 0 1 1
use contact_7  contact_7_50
timestamp 1624857261
transform 1 0 7280 0 1 40253
box 0 0 1 1
use contact_19  contact_19_50
timestamp 1624857261
transform 1 0 7281 0 1 40258
box 0 0 1 1
use and3_dec  and3_dec_25
timestamp 1624857261
transform 1 0 5803 0 1 40290
box 0 -60 2072 490
use contact_17  contact_17_76
timestamp 1624857261
transform 1 0 4904 0 1 40454
box 0 0 1 1
use contact_17  contact_17_75
timestamp 1624857261
transform 1 0 5624 0 1 40544
box 0 0 1 1
use contact_7  contact_7_49
timestamp 1624857261
transform 1 0 6041 0 1 40671
box 0 0 1 1
use contact_19  contact_19_49
timestamp 1624857261
transform 1 0 6042 0 1 40676
box 0 0 1 1
use contact_7  contact_7_328
timestamp 1624857261
transform 1 0 6466 0 1 40671
box 0 0 1 1
use contact_19  contact_19_328
timestamp 1624857261
transform 1 0 6467 0 1 40676
box 0 0 1 1
use contact_7  contact_7_326
timestamp 1624857261
transform 1 0 6898 0 1 40671
box 0 0 1 1
use contact_19  contact_19_326
timestamp 1624857261
transform 1 0 6899 0 1 40676
box 0 0 1 1
use contact_7  contact_7_48
timestamp 1624857261
transform 1 0 7280 0 1 40648
box 0 0 1 1
use contact_19  contact_19_48
timestamp 1624857261
transform 1 0 7281 0 1 40653
box 0 0 1 1
use contact_17  contact_17_73
timestamp 1624857261
transform 1 0 4904 0 1 40858
box 0 0 1 1
use contact_17  contact_17_72
timestamp 1624857261
transform 1 0 5624 0 1 40768
box 0 0 1 1
use and3_dec  and3_dec_24
timestamp 1624857261
transform 1 0 5803 0 -1 41080
box 0 -60 2072 490
use contact_17  contact_17_71
timestamp 1624857261
transform 1 0 4504 0 1 41132
box 0 0 1 1
use contact_17  contact_17_74
timestamp 1624857261
transform 1 0 4744 0 1 40970
box 0 0 1 1
use contact_7  contact_7_47
timestamp 1624857261
transform 1 0 6041 0 1 41087
box 0 0 1 1
use contact_19  contact_19_47
timestamp 1624857261
transform 1 0 6042 0 1 41092
box 0 0 1 1
use contact_7  contact_7_325
timestamp 1624857261
transform 1 0 6466 0 1 41029
box 0 0 1 1
use contact_19  contact_19_325
timestamp 1624857261
transform 1 0 6467 0 1 41034
box 0 0 1 1
use contact_7  contact_7_323
timestamp 1624857261
transform 1 0 6898 0 1 41029
box 0 0 1 1
use contact_19  contact_19_323
timestamp 1624857261
transform 1 0 6899 0 1 41034
box 0 0 1 1
use contact_7  contact_7_46
timestamp 1624857261
transform 1 0 7280 0 1 41043
box 0 0 1 1
use contact_19  contact_19_46
timestamp 1624857261
transform 1 0 7281 0 1 41048
box 0 0 1 1
use contact_17  contact_17_70
timestamp 1624857261
transform 1 0 4984 0 1 41244
box 0 0 1 1
use contact_17  contact_17_69
timestamp 1624857261
transform 1 0 5624 0 1 41334
box 0 0 1 1
use contact_7  contact_7_45
timestamp 1624857261
transform 1 0 6041 0 1 41461
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1624857261
transform 1 0 6042 0 1 41466
box 0 0 1 1
use contact_7  contact_7_322
timestamp 1624857261
transform 1 0 6466 0 1 41461
box 0 0 1 1
use contact_19  contact_19_322
timestamp 1624857261
transform 1 0 6467 0 1 41466
box 0 0 1 1
use contact_7  contact_7_320
timestamp 1624857261
transform 1 0 6898 0 1 41461
box 0 0 1 1
use contact_19  contact_19_320
timestamp 1624857261
transform 1 0 6899 0 1 41466
box 0 0 1 1
use contact_7  contact_7_44
timestamp 1624857261
transform 1 0 7280 0 1 41438
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1624857261
transform 1 0 7281 0 1 41443
box 0 0 1 1
use and3_dec  and3_dec_23
timestamp 1624857261
transform 1 0 5803 0 1 41080
box 0 -60 2072 490
use and3_dec  and3_dec_22
timestamp 1624857261
transform 1 0 5803 0 -1 41870
box 0 -60 2072 490
use contact_17  contact_17_68
timestamp 1624857261
transform 1 0 4584 0 1 41760
box 0 0 1 1
use contact_17  contact_17_67
timestamp 1624857261
transform 1 0 4984 0 1 41648
box 0 0 1 1
use contact_17  contact_17_66
timestamp 1624857261
transform 1 0 5624 0 1 41558
box 0 0 1 1
use contact_17  contact_17_65
timestamp 1624857261
transform 1 0 4664 0 1 41922
box 0 0 1 1
use contact_17  contact_17_64
timestamp 1624857261
transform 1 0 4984 0 1 42034
box 0 0 1 1
use contact_7  contact_7_43
timestamp 1624857261
transform 1 0 6041 0 1 41877
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1624857261
transform 1 0 6042 0 1 41882
box 0 0 1 1
use contact_7  contact_7_319
timestamp 1624857261
transform 1 0 6466 0 1 41819
box 0 0 1 1
use contact_19  contact_19_319
timestamp 1624857261
transform 1 0 6467 0 1 41824
box 0 0 1 1
use contact_7  contact_7_317
timestamp 1624857261
transform 1 0 6898 0 1 41819
box 0 0 1 1
use contact_19  contact_19_317
timestamp 1624857261
transform 1 0 6899 0 1 41824
box 0 0 1 1
use contact_7  contact_7_42
timestamp 1624857261
transform 1 0 7280 0 1 41833
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1624857261
transform 1 0 7281 0 1 41838
box 0 0 1 1
use and3_dec  and3_dec_21
timestamp 1624857261
transform 1 0 5803 0 1 41870
box 0 -60 2072 490
use contact_17  contact_17_63
timestamp 1624857261
transform 1 0 5624 0 1 42124
box 0 0 1 1
use contact_19  contact_19_316
timestamp 1624857261
transform 1 0 6467 0 1 42256
box 0 0 1 1
use contact_7  contact_7_316
timestamp 1624857261
transform 1 0 6466 0 1 42251
box 0 0 1 1
use contact_19  contact_19_314
timestamp 1624857261
transform 1 0 6899 0 1 42256
box 0 0 1 1
use contact_7  contact_7_314
timestamp 1624857261
transform 1 0 6898 0 1 42251
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1624857261
transform 1 0 6042 0 1 42256
box 0 0 1 1
use contact_7  contact_7_41
timestamp 1624857261
transform 1 0 6041 0 1 42251
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1624857261
transform 1 0 7281 0 1 42233
box 0 0 1 1
use contact_7  contact_7_40
timestamp 1624857261
transform 1 0 7280 0 1 42228
box 0 0 1 1
use contact_17  contact_17_62
timestamp 1624857261
transform 1 0 4744 0 1 42550
box 0 0 1 1
use contact_17  contact_17_61
timestamp 1624857261
transform 1 0 4984 0 1 42438
box 0 0 1 1
use contact_17  contact_17_60
timestamp 1624857261
transform 1 0 5624 0 1 42348
box 0 0 1 1
use and3_dec  and3_dec_20
timestamp 1624857261
transform 1 0 5803 0 -1 42660
box 0 -60 2072 490
use contact_7  contact_7_333
timestamp 1624857261
transform 1 0 7676 0 1 39858
box 0 0 1 1
use contact_19  contact_19_333
timestamp 1624857261
transform 1 0 7677 0 1 39863
box 0 0 1 1
use contact_7  contact_7_336
timestamp 1624857261
transform 1 0 7676 0 1 39463
box 0 0 1 1
use contact_19  contact_19_336
timestamp 1624857261
transform 1 0 7677 0 1 39468
box 0 0 1 1
use contact_7  contact_7_324
timestamp 1624857261
transform 1 0 7676 0 1 41043
box 0 0 1 1
use contact_19  contact_19_324
timestamp 1624857261
transform 1 0 7677 0 1 41048
box 0 0 1 1
use contact_7  contact_7_327
timestamp 1624857261
transform 1 0 7676 0 1 40648
box 0 0 1 1
use contact_19  contact_19_327
timestamp 1624857261
transform 1 0 7677 0 1 40653
box 0 0 1 1
use contact_7  contact_7_330
timestamp 1624857261
transform 1 0 7676 0 1 40253
box 0 0 1 1
use contact_19  contact_19_330
timestamp 1624857261
transform 1 0 7677 0 1 40258
box 0 0 1 1
use contact_7  contact_7_318
timestamp 1624857261
transform 1 0 7676 0 1 41833
box 0 0 1 1
use contact_19  contact_19_318
timestamp 1624857261
transform 1 0 7677 0 1 41838
box 0 0 1 1
use contact_7  contact_7_321
timestamp 1624857261
transform 1 0 7676 0 1 41438
box 0 0 1 1
use contact_19  contact_19_321
timestamp 1624857261
transform 1 0 7677 0 1 41443
box 0 0 1 1
use contact_7  contact_7_315
timestamp 1624857261
transform 1 0 7676 0 1 42228
box 0 0 1 1
use contact_19  contact_19_315
timestamp 1624857261
transform 1 0 7677 0 1 42233
box 0 0 1 1
use contact_17  contact_17_59
timestamp 1624857261
transform 1 0 4504 0 1 42712
box 0 0 1 1
use contact_17  contact_17_58
timestamp 1624857261
transform 1 0 5064 0 1 42824
box 0 0 1 1
use contact_7  contact_7_39
timestamp 1624857261
transform 1 0 6041 0 1 42667
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1624857261
transform 1 0 6042 0 1 42672
box 0 0 1 1
use contact_7  contact_7_313
timestamp 1624857261
transform 1 0 6466 0 1 42609
box 0 0 1 1
use contact_19  contact_19_313
timestamp 1624857261
transform 1 0 6467 0 1 42614
box 0 0 1 1
use contact_7  contact_7_311
timestamp 1624857261
transform 1 0 6898 0 1 42609
box 0 0 1 1
use contact_19  contact_19_311
timestamp 1624857261
transform 1 0 6899 0 1 42614
box 0 0 1 1
use contact_7  contact_7_38
timestamp 1624857261
transform 1 0 7280 0 1 42623
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1624857261
transform 1 0 7281 0 1 42628
box 0 0 1 1
use contact_17  contact_17_54
timestamp 1624857261
transform 1 0 5624 0 1 43138
box 0 0 1 1
use contact_17  contact_17_57
timestamp 1624857261
transform 1 0 5624 0 1 42914
box 0 0 1 1
use contact_7  contact_7_37
timestamp 1624857261
transform 1 0 6041 0 1 43041
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1624857261
transform 1 0 6042 0 1 43046
box 0 0 1 1
use contact_7  contact_7_310
timestamp 1624857261
transform 1 0 6466 0 1 43041
box 0 0 1 1
use contact_19  contact_19_310
timestamp 1624857261
transform 1 0 6467 0 1 43046
box 0 0 1 1
use contact_7  contact_7_308
timestamp 1624857261
transform 1 0 6898 0 1 43041
box 0 0 1 1
use contact_19  contact_19_308
timestamp 1624857261
transform 1 0 6899 0 1 43046
box 0 0 1 1
use contact_7  contact_7_36
timestamp 1624857261
transform 1 0 7280 0 1 43018
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1624857261
transform 1 0 7281 0 1 43023
box 0 0 1 1
use and3_dec  and3_dec_19
timestamp 1624857261
transform 1 0 5803 0 1 42660
box 0 -60 2072 490
use and3_dec  and3_dec_18
timestamp 1624857261
transform 1 0 5803 0 -1 43450
box 0 -60 2072 490
use contact_17  contact_17_56
timestamp 1624857261
transform 1 0 4584 0 1 43340
box 0 0 1 1
use contact_17  contact_17_55
timestamp 1624857261
transform 1 0 5064 0 1 43228
box 0 0 1 1
use contact_19  contact_19_307
timestamp 1624857261
transform 1 0 6467 0 1 43404
box 0 0 1 1
use contact_7  contact_7_307
timestamp 1624857261
transform 1 0 6466 0 1 43399
box 0 0 1 1
use contact_19  contact_19_305
timestamp 1624857261
transform 1 0 6899 0 1 43404
box 0 0 1 1
use contact_7  contact_7_305
timestamp 1624857261
transform 1 0 6898 0 1 43399
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1624857261
transform 1 0 7281 0 1 43418
box 0 0 1 1
use contact_7  contact_7_34
timestamp 1624857261
transform 1 0 7280 0 1 43413
box 0 0 1 1
use contact_17  contact_17_53
timestamp 1624857261
transform 1 0 4664 0 1 43502
box 0 0 1 1
use contact_17  contact_17_52
timestamp 1624857261
transform 1 0 5064 0 1 43614
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1624857261
transform 1 0 6042 0 1 43462
box 0 0 1 1
use contact_7  contact_7_35
timestamp 1624857261
transform 1 0 6041 0 1 43457
box 0 0 1 1
use and3_dec  and3_dec_17
timestamp 1624857261
transform 1 0 5803 0 1 43450
box 0 -60 2072 490
use contact_17  contact_17_48
timestamp 1624857261
transform 1 0 5624 0 1 43928
box 0 0 1 1
use contact_17  contact_17_51
timestamp 1624857261
transform 1 0 5624 0 1 43704
box 0 0 1 1
use contact_7  contact_7_33
timestamp 1624857261
transform 1 0 6041 0 1 43831
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1624857261
transform 1 0 6042 0 1 43836
box 0 0 1 1
use contact_7  contact_7_304
timestamp 1624857261
transform 1 0 6466 0 1 43831
box 0 0 1 1
use contact_19  contact_19_304
timestamp 1624857261
transform 1 0 6467 0 1 43836
box 0 0 1 1
use contact_7  contact_7_302
timestamp 1624857261
transform 1 0 6898 0 1 43831
box 0 0 1 1
use contact_19  contact_19_302
timestamp 1624857261
transform 1 0 6899 0 1 43836
box 0 0 1 1
use contact_7  contact_7_32
timestamp 1624857261
transform 1 0 7280 0 1 43808
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1624857261
transform 1 0 7281 0 1 43813
box 0 0 1 1
use contact_17  contact_17_50
timestamp 1624857261
transform 1 0 4744 0 1 44130
box 0 0 1 1
use contact_17  contact_17_49
timestamp 1624857261
transform 1 0 5064 0 1 44018
box 0 0 1 1
use contact_19  contact_19_301
timestamp 1624857261
transform 1 0 6467 0 1 44194
box 0 0 1 1
use contact_7  contact_7_301
timestamp 1624857261
transform 1 0 6466 0 1 44189
box 0 0 1 1
use contact_19  contact_19_299
timestamp 1624857261
transform 1 0 6899 0 1 44194
box 0 0 1 1
use contact_7  contact_7_299
timestamp 1624857261
transform 1 0 6898 0 1 44189
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1624857261
transform 1 0 7281 0 1 44208
box 0 0 1 1
use contact_7  contact_7_30
timestamp 1624857261
transform 1 0 7280 0 1 44203
box 0 0 1 1
use and3_dec  and3_dec_16
timestamp 1624857261
transform 1 0 5803 0 -1 44240
box 0 -60 2072 490
use and3_dec  and3_dec_15
timestamp 1624857261
transform 1 0 5803 0 1 44240
box 0 -60 2072 490
use contact_17  contact_17_47
timestamp 1624857261
transform 1 0 4504 0 1 44292
box 0 0 1 1
use contact_17  contact_17_46
timestamp 1624857261
transform 1 0 4824 0 1 44404
box 0 0 1 1
use contact_17  contact_17_45
timestamp 1624857261
transform 1 0 5704 0 1 44494
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1624857261
transform 1 0 6042 0 1 44252
box 0 0 1 1
use contact_7  contact_7_31
timestamp 1624857261
transform 1 0 6041 0 1 44247
box 0 0 1 1
use contact_17  contact_17_42
timestamp 1624857261
transform 1 0 5704 0 1 44718
box 0 0 1 1
use contact_19  contact_19_298
timestamp 1624857261
transform 1 0 6467 0 1 44626
box 0 0 1 1
use contact_7  contact_7_298
timestamp 1624857261
transform 1 0 6466 0 1 44621
box 0 0 1 1
use contact_19  contact_19_296
timestamp 1624857261
transform 1 0 6899 0 1 44626
box 0 0 1 1
use contact_7  contact_7_296
timestamp 1624857261
transform 1 0 6898 0 1 44621
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1624857261
transform 1 0 6042 0 1 44626
box 0 0 1 1
use contact_7  contact_7_29
timestamp 1624857261
transform 1 0 6041 0 1 44621
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1624857261
transform 1 0 7281 0 1 44603
box 0 0 1 1
use contact_7  contact_7_28
timestamp 1624857261
transform 1 0 7280 0 1 44598
box 0 0 1 1
use and3_dec  and3_dec_14
timestamp 1624857261
transform 1 0 5803 0 -1 45030
box 0 -60 2072 490
use contact_17  contact_17_43
timestamp 1624857261
transform 1 0 4824 0 1 44808
box 0 0 1 1
use contact_17  contact_17_44
timestamp 1624857261
transform 1 0 4584 0 1 44920
box 0 0 1 1
use contact_7  contact_7_27
timestamp 1624857261
transform 1 0 6041 0 1 45037
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1624857261
transform 1 0 6042 0 1 45042
box 0 0 1 1
use contact_7  contact_7_295
timestamp 1624857261
transform 1 0 6466 0 1 44979
box 0 0 1 1
use contact_19  contact_19_295
timestamp 1624857261
transform 1 0 6467 0 1 44984
box 0 0 1 1
use contact_7  contact_7_293
timestamp 1624857261
transform 1 0 6898 0 1 44979
box 0 0 1 1
use contact_19  contact_19_293
timestamp 1624857261
transform 1 0 6899 0 1 44984
box 0 0 1 1
use contact_7  contact_7_26
timestamp 1624857261
transform 1 0 7280 0 1 44993
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1624857261
transform 1 0 7281 0 1 44998
box 0 0 1 1
use contact_17  contact_17_41
timestamp 1624857261
transform 1 0 4664 0 1 45082
box 0 0 1 1
use contact_17  contact_17_40
timestamp 1624857261
transform 1 0 4824 0 1 45194
box 0 0 1 1
use contact_17  contact_17_39
timestamp 1624857261
transform 1 0 5704 0 1 45284
box 0 0 1 1
use and3_dec  and3_dec_13
timestamp 1624857261
transform 1 0 5803 0 1 45030
box 0 -60 2072 490
use and3_dec  and3_dec_12
timestamp 1624857261
transform 1 0 5803 0 -1 45820
box 0 -60 2072 490
use contact_17  contact_17_37
timestamp 1624857261
transform 1 0 4824 0 1 45598
box 0 0 1 1
use contact_7  contact_7_25
timestamp 1624857261
transform 1 0 6041 0 1 45411
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1624857261
transform 1 0 6042 0 1 45416
box 0 0 1 1
use contact_17  contact_17_36
timestamp 1624857261
transform 1 0 5704 0 1 45508
box 0 0 1 1
use contact_7  contact_7_292
timestamp 1624857261
transform 1 0 6466 0 1 45411
box 0 0 1 1
use contact_19  contact_19_292
timestamp 1624857261
transform 1 0 6467 0 1 45416
box 0 0 1 1
use contact_7  contact_7_290
timestamp 1624857261
transform 1 0 6898 0 1 45411
box 0 0 1 1
use contact_19  contact_19_290
timestamp 1624857261
transform 1 0 6899 0 1 45416
box 0 0 1 1
use contact_7  contact_7_24
timestamp 1624857261
transform 1 0 7280 0 1 45388
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1624857261
transform 1 0 7281 0 1 45393
box 0 0 1 1
use contact_17  contact_17_35
timestamp 1624857261
transform 1 0 4504 0 1 45872
box 0 0 1 1
use contact_17  contact_17_38
timestamp 1624857261
transform 1 0 4744 0 1 45710
box 0 0 1 1
use contact_7  contact_7_23
timestamp 1624857261
transform 1 0 6041 0 1 45827
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1624857261
transform 1 0 6042 0 1 45832
box 0 0 1 1
use contact_7  contact_7_289
timestamp 1624857261
transform 1 0 6466 0 1 45769
box 0 0 1 1
use contact_19  contact_19_289
timestamp 1624857261
transform 1 0 6467 0 1 45774
box 0 0 1 1
use contact_7  contact_7_287
timestamp 1624857261
transform 1 0 6898 0 1 45769
box 0 0 1 1
use contact_19  contact_19_287
timestamp 1624857261
transform 1 0 6899 0 1 45774
box 0 0 1 1
use contact_7  contact_7_22
timestamp 1624857261
transform 1 0 7280 0 1 45783
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1624857261
transform 1 0 7281 0 1 45788
box 0 0 1 1
use and3_dec  and3_dec_11
timestamp 1624857261
transform 1 0 5803 0 1 45820
box 0 -60 2072 490
use contact_7  contact_7_306
timestamp 1624857261
transform 1 0 7676 0 1 43413
box 0 0 1 1
use contact_19  contact_19_306
timestamp 1624857261
transform 1 0 7677 0 1 43418
box 0 0 1 1
use contact_7  contact_7_309
timestamp 1624857261
transform 1 0 7676 0 1 43018
box 0 0 1 1
use contact_19  contact_19_309
timestamp 1624857261
transform 1 0 7677 0 1 43023
box 0 0 1 1
use contact_7  contact_7_312
timestamp 1624857261
transform 1 0 7676 0 1 42623
box 0 0 1 1
use contact_19  contact_19_312
timestamp 1624857261
transform 1 0 7677 0 1 42628
box 0 0 1 1
use contact_7  contact_7_300
timestamp 1624857261
transform 1 0 7676 0 1 44203
box 0 0 1 1
use contact_19  contact_19_300
timestamp 1624857261
transform 1 0 7677 0 1 44208
box 0 0 1 1
use contact_7  contact_7_303
timestamp 1624857261
transform 1 0 7676 0 1 43808
box 0 0 1 1
use contact_19  contact_19_303
timestamp 1624857261
transform 1 0 7677 0 1 43813
box 0 0 1 1
use contact_7  contact_7_294
timestamp 1624857261
transform 1 0 7676 0 1 44993
box 0 0 1 1
use contact_19  contact_19_294
timestamp 1624857261
transform 1 0 7677 0 1 44998
box 0 0 1 1
use contact_7  contact_7_297
timestamp 1624857261
transform 1 0 7676 0 1 44598
box 0 0 1 1
use contact_19  contact_19_297
timestamp 1624857261
transform 1 0 7677 0 1 44603
box 0 0 1 1
use contact_7  contact_7_288
timestamp 1624857261
transform 1 0 7676 0 1 45783
box 0 0 1 1
use contact_19  contact_19_288
timestamp 1624857261
transform 1 0 7677 0 1 45788
box 0 0 1 1
use contact_7  contact_7_291
timestamp 1624857261
transform 1 0 7676 0 1 45388
box 0 0 1 1
use contact_19  contact_19_291
timestamp 1624857261
transform 1 0 7677 0 1 45393
box 0 0 1 1
use contact_17  contact_17_34
timestamp 1624857261
transform 1 0 4904 0 1 45984
box 0 0 1 1
use contact_17  contact_17_33
timestamp 1624857261
transform 1 0 5704 0 1 46074
box 0 0 1 1
use contact_17  contact_17_31
timestamp 1624857261
transform 1 0 4904 0 1 46388
box 0 0 1 1
use contact_7  contact_7_21
timestamp 1624857261
transform 1 0 6041 0 1 46201
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1624857261
transform 1 0 6042 0 1 46206
box 0 0 1 1
use contact_17  contact_17_30
timestamp 1624857261
transform 1 0 5704 0 1 46298
box 0 0 1 1
use contact_7  contact_7_286
timestamp 1624857261
transform 1 0 6466 0 1 46201
box 0 0 1 1
use contact_19  contact_19_286
timestamp 1624857261
transform 1 0 6467 0 1 46206
box 0 0 1 1
use contact_7  contact_7_284
timestamp 1624857261
transform 1 0 6898 0 1 46201
box 0 0 1 1
use contact_19  contact_19_284
timestamp 1624857261
transform 1 0 6899 0 1 46206
box 0 0 1 1
use contact_7  contact_7_20
timestamp 1624857261
transform 1 0 7280 0 1 46178
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1624857261
transform 1 0 7281 0 1 46183
box 0 0 1 1
use and3_dec  and3_dec_10
timestamp 1624857261
transform 1 0 5803 0 -1 46610
box 0 -60 2072 490
use contact_17  contact_17_29
timestamp 1624857261
transform 1 0 4664 0 1 46662
box 0 0 1 1
use contact_17  contact_17_32
timestamp 1624857261
transform 1 0 4584 0 1 46500
box 0 0 1 1
use contact_7  contact_7_19
timestamp 1624857261
transform 1 0 6041 0 1 46617
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1624857261
transform 1 0 6042 0 1 46622
box 0 0 1 1
use contact_7  contact_7_283
timestamp 1624857261
transform 1 0 6466 0 1 46559
box 0 0 1 1
use contact_19  contact_19_283
timestamp 1624857261
transform 1 0 6467 0 1 46564
box 0 0 1 1
use contact_7  contact_7_281
timestamp 1624857261
transform 1 0 6898 0 1 46559
box 0 0 1 1
use contact_19  contact_19_281
timestamp 1624857261
transform 1 0 6899 0 1 46564
box 0 0 1 1
use contact_7  contact_7_18
timestamp 1624857261
transform 1 0 7280 0 1 46573
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1624857261
transform 1 0 7281 0 1 46578
box 0 0 1 1
use contact_17  contact_17_28
timestamp 1624857261
transform 1 0 4904 0 1 46774
box 0 0 1 1
use contact_17  contact_17_27
timestamp 1624857261
transform 1 0 5704 0 1 46864
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1624857261
transform 1 0 7281 0 1 46973
box 0 0 1 1
use contact_7  contact_7_16
timestamp 1624857261
transform 1 0 7280 0 1 46968
box 0 0 1 1
use and3_dec  and3_dec_9
timestamp 1624857261
transform 1 0 5803 0 1 46610
box 0 -60 2072 490
use and3_dec  and3_dec_8
timestamp 1624857261
transform 1 0 5803 0 -1 47400
box 0 -60 2072 490
use contact_17  contact_17_25
timestamp 1624857261
transform 1 0 4904 0 1 47178
box 0 0 1 1
use contact_17  contact_17_24
timestamp 1624857261
transform 1 0 5704 0 1 47088
box 0 0 1 1
use contact_19  contact_19_280
timestamp 1624857261
transform 1 0 6467 0 1 46996
box 0 0 1 1
use contact_7  contact_7_280
timestamp 1624857261
transform 1 0 6466 0 1 46991
box 0 0 1 1
use contact_19  contact_19_278
timestamp 1624857261
transform 1 0 6899 0 1 46996
box 0 0 1 1
use contact_7  contact_7_278
timestamp 1624857261
transform 1 0 6898 0 1 46991
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1624857261
transform 1 0 6042 0 1 46996
box 0 0 1 1
use contact_7  contact_7_17
timestamp 1624857261
transform 1 0 6041 0 1 46991
box 0 0 1 1
use contact_17  contact_17_23
timestamp 1624857261
transform 1 0 4504 0 1 47452
box 0 0 1 1
use contact_17  contact_17_26
timestamp 1624857261
transform 1 0 4744 0 1 47290
box 0 0 1 1
use contact_7  contact_7_15
timestamp 1624857261
transform 1 0 6041 0 1 47407
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1624857261
transform 1 0 6042 0 1 47412
box 0 0 1 1
use contact_7  contact_7_277
timestamp 1624857261
transform 1 0 6466 0 1 47349
box 0 0 1 1
use contact_19  contact_19_277
timestamp 1624857261
transform 1 0 6467 0 1 47354
box 0 0 1 1
use contact_7  contact_7_275
timestamp 1624857261
transform 1 0 6898 0 1 47349
box 0 0 1 1
use contact_19  contact_19_275
timestamp 1624857261
transform 1 0 6899 0 1 47354
box 0 0 1 1
use contact_7  contact_7_14
timestamp 1624857261
transform 1 0 7280 0 1 47363
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1624857261
transform 1 0 7281 0 1 47368
box 0 0 1 1
use and3_dec  and3_dec_7
timestamp 1624857261
transform 1 0 5803 0 1 47400
box 0 -60 2072 490
use contact_17  contact_17_22
timestamp 1624857261
transform 1 0 4984 0 1 47564
box 0 0 1 1
use contact_7  contact_7_13
timestamp 1624857261
transform 1 0 6041 0 1 47781
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1624857261
transform 1 0 6042 0 1 47786
box 0 0 1 1
use contact_17  contact_17_21
timestamp 1624857261
transform 1 0 5704 0 1 47654
box 0 0 1 1
use contact_7  contact_7_274
timestamp 1624857261
transform 1 0 6466 0 1 47781
box 0 0 1 1
use contact_19  contact_19_274
timestamp 1624857261
transform 1 0 6467 0 1 47786
box 0 0 1 1
use contact_7  contact_7_272
timestamp 1624857261
transform 1 0 6898 0 1 47781
box 0 0 1 1
use contact_19  contact_19_272
timestamp 1624857261
transform 1 0 6899 0 1 47786
box 0 0 1 1
use contact_7  contact_7_12
timestamp 1624857261
transform 1 0 7280 0 1 47758
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1624857261
transform 1 0 7281 0 1 47763
box 0 0 1 1
use contact_17  contact_17_19
timestamp 1624857261
transform 1 0 4984 0 1 47968
box 0 0 1 1
use contact_17  contact_17_18
timestamp 1624857261
transform 1 0 5704 0 1 47878
box 0 0 1 1
use and3_dec  and3_dec_6
timestamp 1624857261
transform 1 0 5803 0 -1 48190
box 0 -60 2072 490
use contact_17  contact_17_17
timestamp 1624857261
transform 1 0 4664 0 1 48242
box 0 0 1 1
use contact_17  contact_17_20
timestamp 1624857261
transform 1 0 4584 0 1 48080
box 0 0 1 1
use contact_7  contact_7_11
timestamp 1624857261
transform 1 0 6041 0 1 48197
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1624857261
transform 1 0 6042 0 1 48202
box 0 0 1 1
use contact_7  contact_7_271
timestamp 1624857261
transform 1 0 6466 0 1 48139
box 0 0 1 1
use contact_19  contact_19_271
timestamp 1624857261
transform 1 0 6467 0 1 48144
box 0 0 1 1
use contact_7  contact_7_269
timestamp 1624857261
transform 1 0 6898 0 1 48139
box 0 0 1 1
use contact_19  contact_19_269
timestamp 1624857261
transform 1 0 6899 0 1 48144
box 0 0 1 1
use contact_7  contact_7_10
timestamp 1624857261
transform 1 0 7280 0 1 48153
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1624857261
transform 1 0 7281 0 1 48158
box 0 0 1 1
use contact_17  contact_17_16
timestamp 1624857261
transform 1 0 4984 0 1 48354
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1624857261
transform 1 0 6041 0 1 48571
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1624857261
transform 1 0 6042 0 1 48576
box 0 0 1 1
use contact_17  contact_17_15
timestamp 1624857261
transform 1 0 5704 0 1 48444
box 0 0 1 1
use contact_7  contact_7_268
timestamp 1624857261
transform 1 0 6466 0 1 48571
box 0 0 1 1
use contact_19  contact_19_268
timestamp 1624857261
transform 1 0 6467 0 1 48576
box 0 0 1 1
use contact_7  contact_7_266
timestamp 1624857261
transform 1 0 6898 0 1 48571
box 0 0 1 1
use contact_19  contact_19_266
timestamp 1624857261
transform 1 0 6899 0 1 48576
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1624857261
transform 1 0 7280 0 1 48548
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1624857261
transform 1 0 7281 0 1 48553
box 0 0 1 1
use and3_dec  and3_dec_5
timestamp 1624857261
transform 1 0 5803 0 1 48190
box 0 -60 2072 490
use and3_dec  and3_dec_4
timestamp 1624857261
transform 1 0 5803 0 -1 48980
box 0 -60 2072 490
use contact_17  contact_17_14
timestamp 1624857261
transform 1 0 4744 0 1 48870
box 0 0 1 1
use contact_17  contact_17_13
timestamp 1624857261
transform 1 0 4984 0 1 48758
box 0 0 1 1
use contact_17  contact_17_12
timestamp 1624857261
transform 1 0 5704 0 1 48668
box 0 0 1 1
use contact_17  contact_17_11
timestamp 1624857261
transform 1 0 4504 0 1 49032
box 0 0 1 1
use contact_17  contact_17_10
timestamp 1624857261
transform 1 0 5064 0 1 49144
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1624857261
transform 1 0 6041 0 1 48987
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1624857261
transform 1 0 6042 0 1 48992
box 0 0 1 1
use contact_7  contact_7_265
timestamp 1624857261
transform 1 0 6466 0 1 48929
box 0 0 1 1
use contact_19  contact_19_265
timestamp 1624857261
transform 1 0 6467 0 1 48934
box 0 0 1 1
use contact_7  contact_7_263
timestamp 1624857261
transform 1 0 6898 0 1 48929
box 0 0 1 1
use contact_19  contact_19_263
timestamp 1624857261
transform 1 0 6899 0 1 48934
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1624857261
transform 1 0 7280 0 1 48943
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1624857261
transform 1 0 7281 0 1 48948
box 0 0 1 1
use and3_dec  and3_dec_3
timestamp 1624857261
transform 1 0 5803 0 1 48980
box 0 -60 2072 490
use contact_7  contact_7_282
timestamp 1624857261
transform 1 0 7676 0 1 46573
box 0 0 1 1
use contact_19  contact_19_282
timestamp 1624857261
transform 1 0 7677 0 1 46578
box 0 0 1 1
use contact_7  contact_7_285
timestamp 1624857261
transform 1 0 7676 0 1 46178
box 0 0 1 1
use contact_19  contact_19_285
timestamp 1624857261
transform 1 0 7677 0 1 46183
box 0 0 1 1
use contact_7  contact_7_276
timestamp 1624857261
transform 1 0 7676 0 1 47363
box 0 0 1 1
use contact_19  contact_19_276
timestamp 1624857261
transform 1 0 7677 0 1 47368
box 0 0 1 1
use contact_7  contact_7_279
timestamp 1624857261
transform 1 0 7676 0 1 46968
box 0 0 1 1
use contact_19  contact_19_279
timestamp 1624857261
transform 1 0 7677 0 1 46973
box 0 0 1 1
use contact_7  contact_7_270
timestamp 1624857261
transform 1 0 7676 0 1 48153
box 0 0 1 1
use contact_19  contact_19_270
timestamp 1624857261
transform 1 0 7677 0 1 48158
box 0 0 1 1
use contact_7  contact_7_273
timestamp 1624857261
transform 1 0 7676 0 1 47758
box 0 0 1 1
use contact_19  contact_19_273
timestamp 1624857261
transform 1 0 7677 0 1 47763
box 0 0 1 1
use contact_7  contact_7_264
timestamp 1624857261
transform 1 0 7676 0 1 48943
box 0 0 1 1
use contact_19  contact_19_264
timestamp 1624857261
transform 1 0 7677 0 1 48948
box 0 0 1 1
use contact_7  contact_7_267
timestamp 1624857261
transform 1 0 7676 0 1 48548
box 0 0 1 1
use contact_19  contact_19_267
timestamp 1624857261
transform 1 0 7677 0 1 48553
box 0 0 1 1
use contact_17  contact_17_9
timestamp 1624857261
transform 1 0 5704 0 1 49234
box 0 0 1 1
use contact_19  contact_19_262
timestamp 1624857261
transform 1 0 6467 0 1 49366
box 0 0 1 1
use contact_7  contact_7_262
timestamp 1624857261
transform 1 0 6466 0 1 49361
box 0 0 1 1
use contact_19  contact_19_260
timestamp 1624857261
transform 1 0 6899 0 1 49366
box 0 0 1 1
use contact_7  contact_7_260
timestamp 1624857261
transform 1 0 6898 0 1 49361
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1624857261
transform 1 0 6042 0 1 49366
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1624857261
transform 1 0 6041 0 1 49361
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1624857261
transform 1 0 7281 0 1 49343
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1624857261
transform 1 0 7280 0 1 49338
box 0 0 1 1
use contact_17  contact_17_8
timestamp 1624857261
transform 1 0 4584 0 1 49660
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1624857261
transform 1 0 5064 0 1 49548
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1624857261
transform 1 0 5704 0 1 49458
box 0 0 1 1
use and3_dec  and3_dec_2
timestamp 1624857261
transform 1 0 5803 0 -1 49770
box 0 -60 2072 490
use contact_17  contact_17_5
timestamp 1624857261
transform 1 0 4664 0 1 49822
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1624857261
transform 1 0 5064 0 1 49934
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1624857261
transform 1 0 6041 0 1 49777
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1624857261
transform 1 0 6042 0 1 49782
box 0 0 1 1
use contact_7  contact_7_259
timestamp 1624857261
transform 1 0 6466 0 1 49719
box 0 0 1 1
use contact_19  contact_19_259
timestamp 1624857261
transform 1 0 6467 0 1 49724
box 0 0 1 1
use contact_7  contact_7_257
timestamp 1624857261
transform 1 0 6898 0 1 49719
box 0 0 1 1
use contact_19  contact_19_257
timestamp 1624857261
transform 1 0 6899 0 1 49724
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1624857261
transform 1 0 7280 0 1 49733
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1624857261
transform 1 0 7281 0 1 49738
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1624857261
transform 1 0 6041 0 1 50151
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1624857261
transform 1 0 6042 0 1 50156
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1624857261
transform 1 0 5704 0 1 50248
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1624857261
transform 1 0 5704 0 1 50024
box 0 0 1 1
use contact_7  contact_7_256
timestamp 1624857261
transform 1 0 6466 0 1 50151
box 0 0 1 1
use contact_19  contact_19_256
timestamp 1624857261
transform 1 0 6467 0 1 50156
box 0 0 1 1
use contact_7  contact_7_254
timestamp 1624857261
transform 1 0 6898 0 1 50151
box 0 0 1 1
use contact_19  contact_19_254
timestamp 1624857261
transform 1 0 6899 0 1 50156
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1624857261
transform 1 0 7280 0 1 50128
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1624857261
transform 1 0 7281 0 1 50133
box 0 0 1 1
use and3_dec  and3_dec_1
timestamp 1624857261
transform 1 0 5803 0 1 49770
box 0 -60 2072 490
use and3_dec  and3_dec_0
timestamp 1624857261
transform 1 0 5803 0 -1 50560
box 0 -60 2072 490
use contact_17  contact_17_1
timestamp 1624857261
transform 1 0 5064 0 1 50338
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1624857261
transform 1 0 4744 0 1 50450
box 0 0 1 1
use contact_19  contact_19_261
timestamp 1624857261
transform 1 0 7677 0 1 49343
box 0 0 1 1
use contact_7  contact_7_261
timestamp 1624857261
transform 1 0 7676 0 1 49338
box 0 0 1 1
use contact_19  contact_19_258
timestamp 1624857261
transform 1 0 7677 0 1 49738
box 0 0 1 1
use contact_7  contact_7_258
timestamp 1624857261
transform 1 0 7676 0 1 49733
box 0 0 1 1
use contact_19  contact_19_255
timestamp 1624857261
transform 1 0 7677 0 1 50133
box 0 0 1 1
use contact_7  contact_7_255
timestamp 1624857261
transform 1 0 7676 0 1 50128
box 0 0 1 1
<< labels >>
rlabel metal1 s 19 0 47 7900 4 addr_0
port 1 se
rlabel metal1 s 99 0 127 7900 4 addr_1
port 2 se
rlabel metal1 s 179 0 207 7900 4 addr_2
port 3 se
rlabel metal1 s 259 0 287 7900 4 addr_3
port 4 se
rlabel metal1 s 339 0 367 7900 4 addr_4
port 5 se
rlabel metal1 s 419 0 447 7900 4 addr_5
port 6 se
rlabel metal1 s 499 0 527 7900 4 addr_6
port 7 se
rlabel locali s 7568 120 7568 120 4 decode_0
port 8 se
rlabel locali s 7568 670 7568 670 4 decode_1
port 9 se
rlabel locali s 7568 910 7568 910 4 decode_2
port 10 se
rlabel locali s 7568 1460 7568 1460 4 decode_3
port 11 se
rlabel locali s 7568 1700 7568 1700 4 decode_4
port 12 se
rlabel locali s 7568 2250 7568 2250 4 decode_5
port 13 se
rlabel locali s 7568 2490 7568 2490 4 decode_6
port 14 se
rlabel locali s 7568 3040 7568 3040 4 decode_7
port 15 se
rlabel locali s 7568 3280 7568 3280 4 decode_8
port 16 se
rlabel locali s 7568 3830 7568 3830 4 decode_9
port 17 se
rlabel locali s 7568 4070 7568 4070 4 decode_10
port 18 se
rlabel locali s 7568 4620 7568 4620 4 decode_11
port 19 se
rlabel locali s 7568 4860 7568 4860 4 decode_12
port 20 se
rlabel locali s 7568 5410 7568 5410 4 decode_13
port 21 se
rlabel locali s 7568 5650 7568 5650 4 decode_14
port 22 se
rlabel locali s 7568 6200 7568 6200 4 decode_15
port 23 se
rlabel locali s 7568 6440 7568 6440 4 decode_16
port 24 se
rlabel locali s 7568 6990 7568 6990 4 decode_17
port 25 se
rlabel locali s 7568 7230 7568 7230 4 decode_18
port 26 se
rlabel locali s 7568 7780 7568 7780 4 decode_19
port 27 se
rlabel locali s 7568 8020 7568 8020 4 decode_20
port 28 se
rlabel locali s 7568 8570 7568 8570 4 decode_21
port 29 se
rlabel locali s 7568 8810 7568 8810 4 decode_22
port 30 se
rlabel locali s 7568 9360 7568 9360 4 decode_23
port 31 se
rlabel locali s 7568 9600 7568 9600 4 decode_24
port 32 se
rlabel locali s 7568 10150 7568 10150 4 decode_25
port 33 se
rlabel locali s 7568 10390 7568 10390 4 decode_26
port 34 se
rlabel locali s 7568 10940 7568 10940 4 decode_27
port 35 se
rlabel locali s 7568 11180 7568 11180 4 decode_28
port 36 se
rlabel locali s 7568 11730 7568 11730 4 decode_29
port 37 se
rlabel locali s 7568 11970 7568 11970 4 decode_30
port 38 se
rlabel locali s 7568 12520 7568 12520 4 decode_31
port 39 se
rlabel locali s 7568 12760 7568 12760 4 decode_32
port 40 se
rlabel locali s 7568 13310 7568 13310 4 decode_33
port 41 se
rlabel locali s 7568 13550 7568 13550 4 decode_34
port 42 se
rlabel locali s 7568 14100 7568 14100 4 decode_35
port 43 se
rlabel locali s 7568 14340 7568 14340 4 decode_36
port 44 se
rlabel locali s 7568 14890 7568 14890 4 decode_37
port 45 se
rlabel locali s 7568 15130 7568 15130 4 decode_38
port 46 se
rlabel locali s 7568 15680 7568 15680 4 decode_39
port 47 se
rlabel locali s 7568 15920 7568 15920 4 decode_40
port 48 se
rlabel locali s 7568 16470 7568 16470 4 decode_41
port 49 se
rlabel locali s 7568 16710 7568 16710 4 decode_42
port 50 se
rlabel locali s 7568 17260 7568 17260 4 decode_43
port 51 se
rlabel locali s 7568 17500 7568 17500 4 decode_44
port 52 se
rlabel locali s 7568 18050 7568 18050 4 decode_45
port 53 se
rlabel locali s 7568 18290 7568 18290 4 decode_46
port 54 se
rlabel locali s 7568 18840 7568 18840 4 decode_47
port 55 se
rlabel locali s 7568 19080 7568 19080 4 decode_48
port 56 se
rlabel locali s 7568 19630 7568 19630 4 decode_49
port 57 se
rlabel locali s 7568 19870 7568 19870 4 decode_50
port 58 se
rlabel locali s 7568 20420 7568 20420 4 decode_51
port 59 se
rlabel locali s 7568 20660 7568 20660 4 decode_52
port 60 se
rlabel locali s 7568 21210 7568 21210 4 decode_53
port 61 se
rlabel locali s 7568 21450 7568 21450 4 decode_54
port 62 se
rlabel locali s 7568 22000 7568 22000 4 decode_55
port 63 se
rlabel locali s 7568 22240 7568 22240 4 decode_56
port 64 se
rlabel locali s 7568 22790 7568 22790 4 decode_57
port 65 se
rlabel locali s 7568 23030 7568 23030 4 decode_58
port 66 se
rlabel locali s 7568 23580 7568 23580 4 decode_59
port 67 se
rlabel locali s 7568 23820 7568 23820 4 decode_60
port 68 se
rlabel locali s 7568 24370 7568 24370 4 decode_61
port 69 se
rlabel locali s 7568 24610 7568 24610 4 decode_62
port 70 se
rlabel locali s 7568 25160 7568 25160 4 decode_63
port 71 se
rlabel locali s 7568 25400 7568 25400 4 decode_64
port 72 se
rlabel locali s 7568 25950 7568 25950 4 decode_65
port 73 se
rlabel locali s 7568 26190 7568 26190 4 decode_66
port 74 se
rlabel locali s 7568 26740 7568 26740 4 decode_67
port 75 se
rlabel locali s 7568 26980 7568 26980 4 decode_68
port 76 se
rlabel locali s 7568 27530 7568 27530 4 decode_69
port 77 se
rlabel locali s 7568 27770 7568 27770 4 decode_70
port 78 se
rlabel locali s 7568 28320 7568 28320 4 decode_71
port 79 se
rlabel locali s 7568 28560 7568 28560 4 decode_72
port 80 se
rlabel locali s 7568 29110 7568 29110 4 decode_73
port 81 se
rlabel locali s 7568 29350 7568 29350 4 decode_74
port 82 se
rlabel locali s 7568 29900 7568 29900 4 decode_75
port 83 se
rlabel locali s 7568 30140 7568 30140 4 decode_76
port 84 se
rlabel locali s 7568 30690 7568 30690 4 decode_77
port 85 se
rlabel locali s 7568 30930 7568 30930 4 decode_78
port 86 se
rlabel locali s 7568 31480 7568 31480 4 decode_79
port 87 se
rlabel locali s 7568 31720 7568 31720 4 decode_80
port 88 se
rlabel locali s 7568 32270 7568 32270 4 decode_81
port 89 se
rlabel locali s 7568 32510 7568 32510 4 decode_82
port 90 se
rlabel locali s 7568 33060 7568 33060 4 decode_83
port 91 se
rlabel locali s 7568 33300 7568 33300 4 decode_84
port 92 se
rlabel locali s 7568 33850 7568 33850 4 decode_85
port 93 se
rlabel locali s 7568 34090 7568 34090 4 decode_86
port 94 se
rlabel locali s 7568 34640 7568 34640 4 decode_87
port 95 se
rlabel locali s 7568 34880 7568 34880 4 decode_88
port 96 se
rlabel locali s 7568 35430 7568 35430 4 decode_89
port 97 se
rlabel locali s 7568 35670 7568 35670 4 decode_90
port 98 se
rlabel locali s 7568 36220 7568 36220 4 decode_91
port 99 se
rlabel locali s 7568 36460 7568 36460 4 decode_92
port 100 se
rlabel locali s 7568 37010 7568 37010 4 decode_93
port 101 se
rlabel locali s 7568 37250 7568 37250 4 decode_94
port 102 se
rlabel locali s 7568 37800 7568 37800 4 decode_95
port 103 se
rlabel locali s 7568 38040 7568 38040 4 decode_96
port 104 se
rlabel locali s 7568 38590 7568 38590 4 decode_97
port 105 se
rlabel locali s 7568 38830 7568 38830 4 decode_98
port 106 se
rlabel locali s 7568 39380 7568 39380 4 decode_99
port 107 se
rlabel locali s 7568 39620 7568 39620 4 decode_100
port 108 se
rlabel locali s 7568 40170 7568 40170 4 decode_101
port 109 se
rlabel locali s 7568 40410 7568 40410 4 decode_102
port 110 se
rlabel locali s 7568 40960 7568 40960 4 decode_103
port 111 se
rlabel locali s 7568 41200 7568 41200 4 decode_104
port 112 se
rlabel locali s 7568 41750 7568 41750 4 decode_105
port 113 se
rlabel locali s 7568 41990 7568 41990 4 decode_106
port 114 se
rlabel locali s 7568 42540 7568 42540 4 decode_107
port 115 se
rlabel locali s 7568 42780 7568 42780 4 decode_108
port 116 se
rlabel locali s 7568 43330 7568 43330 4 decode_109
port 117 se
rlabel locali s 7568 43570 7568 43570 4 decode_110
port 118 se
rlabel locali s 7568 44120 7568 44120 4 decode_111
port 119 se
rlabel locali s 7568 44360 7568 44360 4 decode_112
port 120 se
rlabel locali s 7568 44910 7568 44910 4 decode_113
port 121 se
rlabel locali s 7568 45150 7568 45150 4 decode_114
port 122 se
rlabel locali s 7568 45700 7568 45700 4 decode_115
port 123 se
rlabel locali s 7568 45940 7568 45940 4 decode_116
port 124 se
rlabel locali s 7568 46490 7568 46490 4 decode_117
port 125 se
rlabel locali s 7568 46730 7568 46730 4 decode_118
port 126 se
rlabel locali s 7568 47280 7568 47280 4 decode_119
port 127 se
rlabel locali s 7568 47520 7568 47520 4 decode_120
port 128 se
rlabel locali s 7568 48070 7568 48070 4 decode_121
port 129 se
rlabel locali s 7568 48310 7568 48310 4 decode_122
port 130 se
rlabel locali s 7568 48860 7568 48860 4 decode_123
port 131 se
rlabel locali s 7568 49100 7568 49100 4 decode_124
port 132 se
rlabel locali s 7568 49650 7568 49650 4 decode_125
port 133 se
rlabel locali s 7568 49890 7568 49890 4 decode_126
port 134 se
rlabel locali s 7568 50440 7568 50440 4 decode_127
port 135 se
rlabel metal1 s 4523 0 4551 50588 4 predecode_0
rlabel metal1 s 4603 0 4631 50588 4 predecode_1
rlabel metal1 s 4683 0 4711 50588 4 predecode_2
rlabel metal1 s 4763 0 4791 50588 4 predecode_3
rlabel metal1 s 4843 0 4871 50588 4 predecode_4
rlabel metal1 s 4923 0 4951 50588 4 predecode_5
rlabel metal1 s 5003 0 5031 50588 4 predecode_6
rlabel metal1 s 5083 0 5111 50588 4 predecode_7
rlabel metal1 s 5163 0 5191 50588 4 predecode_8
rlabel metal1 s 5243 0 5271 50588 4 predecode_9
rlabel metal1 s 5323 0 5351 50588 4 predecode_10
rlabel metal1 s 5403 0 5431 50588 4 predecode_11
rlabel metal1 s 5483 0 5511 50588 4 predecode_12
rlabel metal1 s 5563 0 5591 50588 4 predecode_13
rlabel metal1 s 5643 0 5671 50588 4 predecode_14
rlabel metal1 s 5723 0 5751 50588 4 predecode_15
rlabel metal3 s 6450 15737 6548 15835 4 vdd
rlabel metal3 s 6450 4319 6548 4417 4 vdd
rlabel metal3 s 6882 23279 6980 23377 4 vdd
rlabel metal3 s 7660 31551 7758 31649 4 vdd
rlabel metal3 s 6882 22847 6980 22945 4 vdd
rlabel metal3 s 7660 1531 7758 1629 4 vdd
rlabel metal3 s 7660 42611 7758 42709 4 vdd
rlabel metal3 s 6882 14157 6980 14255 4 vdd
rlabel metal3 s 6450 21699 6548 21797 4 vdd
rlabel metal3 s 6450 31537 6548 31635 4 vdd
rlabel metal3 s 6882 2307 6980 2405 4 vdd
rlabel metal3 s 6882 37499 6980 37597 4 vdd
rlabel metal3 s 7660 46561 7758 46659 4 vdd
rlabel metal3 s 6450 5109 6548 5207 4 vdd
rlabel metal3 s 7660 23651 7758 23749 4 vdd
rlabel metal3 s 6882 14947 6980 15045 4 vdd
rlabel metal3 s 3036 5899 3134 5997 4 vdd
rlabel metal3 s 7660 24441 7758 24539 4 vdd
rlabel metal3 s 6450 38289 6548 38387 4 vdd
rlabel metal3 s 7660 46956 7758 47054 4 vdd
rlabel metal3 s 7660 27206 7758 27304 4 vdd
rlabel metal3 s 6882 33907 6980 34005 4 vdd
rlabel metal3 s 7660 26811 7758 26909 4 vdd
rlabel metal3 s 6450 28377 6548 28475 4 vdd
rlabel metal3 s 7660 40636 7758 40734 4 vdd
rlabel metal3 s 7660 2321 7758 2419 4 vdd
rlabel metal3 s 6882 18897 6980 18995 4 vdd
rlabel metal3 s 4246 5876 4344 5974 4 vdd
rlabel metal3 s 7660 27996 7758 28094 4 vdd
rlabel metal3 s 7660 41031 7758 41129 4 vdd
rlabel metal3 s 6882 16169 6980 16267 4 vdd
rlabel metal3 s 7660 32736 7758 32834 4 vdd
rlabel metal3 s 6450 9417 6548 9515 4 vdd
rlabel metal3 s 6882 34339 6980 34437 4 vdd
rlabel metal3 s 6882 32327 6980 32425 4 vdd
rlabel metal3 s 6450 9059 6548 9157 4 vdd
rlabel metal3 s 6450 45757 6548 45855 4 vdd
rlabel metal3 s 7660 45771 7758 45869 4 vdd
rlabel metal3 s 7660 17726 7758 17824 4 vdd
rlabel metal3 s 6882 49707 6980 49805 4 vdd
rlabel metal3 s 7660 14171 7758 14269 4 vdd
rlabel metal3 s 6882 7837 6980 7935 4 vdd
rlabel metal3 s 7660 13381 7758 13479 4 vdd
rlabel metal3 s 6882 17317 6980 17415 4 vdd
rlabel metal3 s 6882 6257 6980 6355 4 vdd
rlabel metal3 s 6450 43819 6548 43917 4 vdd
rlabel metal3 s 6882 1949 6980 2047 4 vdd
rlabel metal3 s 7660 33131 7758 33229 4 vdd
rlabel metal3 s 6882 12577 6980 12675 4 vdd
rlabel metal3 s 7660 11801 7758 11899 4 vdd
rlabel metal3 s 7660 25626 7758 25724 4 vdd
rlabel metal3 s 6882 5467 6980 5565 4 vdd
rlabel metal3 s 7660 19306 7758 19404 4 vdd
rlabel metal3 s 6450 11787 6548 11885 4 vdd
rlabel metal3 s 6450 24427 6548 24525 4 vdd
rlabel metal3 s 6450 46189 6548 46287 4 vdd
rlabel metal3 s 7660 24046 7758 24144 4 vdd
rlabel metal3 s 6450 41807 6548 41905 4 vdd
rlabel metal3 s 4246 346 4344 444 4 vdd
rlabel metal3 s 6450 41449 6548 41547 4 vdd
rlabel metal3 s 6882 7479 6980 7577 4 vdd
rlabel metal3 s 7660 1136 7758 1234 4 vdd
rlabel metal3 s 6882 36709 6980 36807 4 vdd
rlabel metal3 s 6450 45399 6548 45497 4 vdd
rlabel metal3 s 6882 15379 6980 15477 4 vdd
rlabel metal3 s 7660 3506 7758 3604 4 vdd
rlabel metal3 s 6882 38647 6980 38745 4 vdd
rlabel metal3 s 4246 6666 4344 6764 4 vdd
rlabel metal3 s 3471 1143 3569 1241 4 vdd
rlabel metal3 s 3036 6689 3134 6787 4 vdd
rlabel metal3 s 6882 34697 6980 34795 4 vdd
rlabel metal3 s 6882 43029 6980 43127 4 vdd
rlabel metal3 s 6882 47337 6980 47435 4 vdd
rlabel metal3 s 2148 2716 2246 2814 4 vdd
rlabel metal3 s 7660 28786 7758 28884 4 vdd
rlabel metal3 s 6450 727 6548 825 4 vdd
rlabel metal3 s 6882 9849 6980 9947 4 vdd
rlabel metal3 s 7660 44981 7758 45079 4 vdd
rlabel metal3 s 6450 37857 6548 37955 4 vdd
rlabel metal3 s 6450 10207 6548 10305 4 vdd
rlabel metal3 s 6882 19329 6980 19427 4 vdd
rlabel metal3 s 3471 3513 3569 3611 4 vdd
rlabel metal3 s 6450 16527 6548 16625 4 vdd
rlabel metal3 s 6882 45757 6980 45855 4 vdd
rlabel metal3 s 7660 40241 7758 40339 4 vdd
rlabel metal3 s 7660 33526 7758 33624 4 vdd
rlabel metal3 s 6450 7047 6548 7145 4 vdd
rlabel metal3 s 6882 41807 6980 41905 4 vdd
rlabel metal3 s 6450 14157 6548 14255 4 vdd
rlabel metal3 s 6882 18107 6980 18205 4 vdd
rlabel metal3 s 6450 25217 6548 25315 4 vdd
rlabel metal3 s 6882 26797 6980 26895 4 vdd
rlabel metal3 s 6882 43387 6980 43485 4 vdd
rlabel metal3 s 7660 31156 7758 31254 4 vdd
rlabel metal3 s 6882 11787 6980 11885 4 vdd
rlabel metal3 s 6882 27587 6980 27685 4 vdd
rlabel metal3 s 6882 48917 6980 49015 4 vdd
rlabel metal3 s 6882 37857 6980 37955 4 vdd
rlabel metal3 s 7660 346 7758 444 4 vdd
rlabel metal3 s 7660 35896 7758 35994 4 vdd
rlabel metal3 s 6882 21267 6980 21365 4 vdd
rlabel metal3 s 7660 39451 7758 39549 4 vdd
rlabel metal3 s 7660 47351 7758 47449 4 vdd
rlabel metal3 s 6882 17749 6980 17847 4 vdd
rlabel metal3 s 7660 34316 7758 34414 4 vdd
rlabel metal3 s 6450 30747 6548 30845 4 vdd
rlabel metal3 s 7660 1926 7758 2024 4 vdd
rlabel metal3 s 7660 30366 7758 30464 4 vdd
rlabel metal3 s 7660 48141 7758 48239 4 vdd
rlabel metal3 s 6450 5899 6548 5997 4 vdd
rlabel metal3 s 7660 7456 7758 7554 4 vdd
rlabel metal3 s 6882 24859 6980 24957 4 vdd
rlabel metal3 s 7660 11011 7758 11109 4 vdd
rlabel metal3 s 6450 37067 6548 37165 4 vdd
rlabel metal3 s 6450 23637 6548 23735 4 vdd
rlabel metal3 s 6450 26007 6548 26105 4 vdd
rlabel metal3 s 7660 16146 7758 16244 4 vdd
rlabel metal3 s 7660 32341 7758 32439 4 vdd
rlabel metal3 s 1552 5086 1650 5184 4 vdd
rlabel metal3 s 7660 8246 7758 8344 4 vdd
rlabel metal3 s 4246 5086 4344 5184 4 vdd
rlabel metal3 s 6450 50139 6548 50237 4 vdd
rlabel metal3 s 6450 29599 6548 29697 4 vdd
rlabel metal3 s 7660 25231 7758 25329 4 vdd
rlabel metal3 s 6882 37067 6980 37165 4 vdd
rlabel metal3 s 7660 15751 7758 15849 4 vdd
rlabel metal3 s 6882 25649 6980 25747 4 vdd
rlabel metal3 s 6450 5467 6548 5565 4 vdd
rlabel metal3 s 6450 29167 6548 29265 4 vdd
rlabel metal3 s 6450 12577 6548 12675 4 vdd
rlabel metal3 s 6882 46547 6980 46645 4 vdd
rlabel metal3 s 6882 28809 6980 28907 4 vdd
rlabel metal3 s 7660 12986 7758 13084 4 vdd
rlabel metal3 s 7660 20096 7758 20194 4 vdd
rlabel metal3 s 6882 43819 6980 43917 4 vdd
rlabel metal3 s 6882 29957 6980 30055 4 vdd
rlabel metal3 s 7660 27601 7758 27699 4 vdd
rlabel metal3 s 6882 26439 6980 26537 4 vdd
rlabel metal3 s 6882 24427 6980 24525 4 vdd
rlabel metal3 s 6882 4677 6980 4775 4 vdd
rlabel metal3 s 6450 40227 6548 40325 4 vdd
rlabel metal3 s 6450 48127 6548 48225 4 vdd
rlabel metal3 s 6450 33549 6548 33647 4 vdd
rlabel metal3 s 6882 28019 6980 28117 4 vdd
rlabel metal3 s 6450 46547 6548 46645 4 vdd
rlabel metal3 s 6882 20119 6980 20217 4 vdd
rlabel metal3 s 6882 49349 6980 49447 4 vdd
rlabel metal3 s 6450 1159 6548 1257 4 vdd
rlabel metal3 s 6450 1949 6548 2047 4 vdd
rlabel metal3 s 7660 34711 7758 34809 4 vdd
rlabel metal3 s 7660 3901 7758 3999 4 vdd
rlabel metal3 s 6450 8269 6548 8367 4 vdd
rlabel metal3 s 6450 39869 6548 39967 4 vdd
rlabel metal3 s 6450 24859 6548 24957 4 vdd
rlabel metal3 s 7660 9826 7758 9924 4 vdd
rlabel metal3 s 6450 2307 6548 2405 4 vdd
rlabel metal3 s 7660 20491 7758 20589 4 vdd
rlabel metal3 s 7660 16936 7758 17034 4 vdd
rlabel metal3 s 6450 37499 6548 37597 4 vdd
rlabel metal3 s 6450 19329 6548 19427 4 vdd
rlabel metal3 s 7660 24836 7758 24934 4 vdd
rlabel metal3 s 6450 369 6548 467 4 vdd
rlabel metal3 s 7660 22861 7758 22959 4 vdd
rlabel metal3 s 6450 29957 6548 30055 4 vdd
rlabel metal3 s 6450 46979 6548 47077 4 vdd
rlabel metal3 s 7660 36291 7758 36389 4 vdd
rlabel metal3 s 7660 43401 7758 43499 4 vdd
rlabel metal3 s 7660 48931 7758 49029 4 vdd
rlabel metal3 s 6450 22057 6548 22155 4 vdd
rlabel metal3 s 7660 23256 7758 23354 4 vdd
rlabel metal3 s 6450 18107 6548 18205 4 vdd
rlabel metal3 s 6882 39437 6980 39535 4 vdd
rlabel metal3 s 6882 45399 6980 45497 4 vdd
rlabel metal3 s 6450 1517 6548 1615 4 vdd
rlabel metal3 s 6882 18539 6980 18637 4 vdd
rlabel metal3 s 6882 1159 6980 1257 4 vdd
rlabel metal3 s 6450 39079 6548 39177 4 vdd
rlabel metal3 s 6882 15737 6980 15835 4 vdd
rlabel metal3 s 6882 22489 6980 22587 4 vdd
rlabel metal3 s 6882 21699 6980 21797 4 vdd
rlabel metal3 s 7660 28391 7758 28489 4 vdd
rlabel metal3 s 7660 12591 7758 12689 4 vdd
rlabel metal3 s 6450 42597 6548 42695 4 vdd
rlabel metal3 s 6882 5899 6980 5997 4 vdd
rlabel metal3 s 6450 24069 6548 24167 4 vdd
rlabel metal3 s 6882 50139 6980 50237 4 vdd
rlabel metal3 s 6450 16959 6548 17057 4 vdd
rlabel metal3 s 7660 17331 7758 17429 4 vdd
rlabel metal3 s 4246 2716 4344 2814 4 vdd
rlabel metal3 s 7660 47746 7758 47844 4 vdd
rlabel metal3 s 6450 49707 6548 49805 4 vdd
rlabel metal3 s 7660 5086 7758 5184 4 vdd
rlabel metal3 s 3471 353 3569 451 4 vdd
rlabel metal3 s 6882 5109 6980 5207 4 vdd
rlabel metal3 s 6882 35487 6980 35585 4 vdd
rlabel metal3 s 7660 39056 7758 39154 4 vdd
rlabel metal3 s 6450 44177 6548 44275 4 vdd
rlabel metal3 s 6450 28809 6548 28907 4 vdd
rlabel metal3 s 7660 7061 7758 7159 4 vdd
rlabel metal3 s 7660 13776 7758 13874 4 vdd
rlabel metal3 s 6450 22489 6548 22587 4 vdd
rlabel metal3 s 7660 6666 7758 6764 4 vdd
rlabel metal3 s 7660 33921 7758 34019 4 vdd
rlabel metal3 s 6882 41449 6980 41547 4 vdd
rlabel metal3 s 6450 13799 6548 13897 4 vdd
rlabel metal3 s 6450 13367 6548 13465 4 vdd
rlabel metal3 s 7660 42216 7758 42314 4 vdd
rlabel metal3 s 6450 17317 6548 17415 4 vdd
rlabel metal3 s 6450 6689 6548 6787 4 vdd
rlabel metal3 s 7660 21676 7758 21774 4 vdd
rlabel metal3 s 6450 41017 6548 41115 4 vdd
rlabel metal3 s 6882 48559 6980 48657 4 vdd
rlabel metal3 s 6882 2739 6980 2837 4 vdd
rlabel metal3 s 7660 31946 7758 32044 4 vdd
rlabel metal3 s 6882 46189 6980 46287 4 vdd
rlabel metal3 s 6882 31179 6980 31277 4 vdd
rlabel metal3 s 6882 35129 6980 35227 4 vdd
rlabel metal3 s 6450 36277 6548 36375 4 vdd
rlabel metal3 s 6882 9059 6980 9157 4 vdd
rlabel metal3 s 6450 32759 6548 32857 4 vdd
rlabel metal3 s 6882 26007 6980 26105 4 vdd
rlabel metal3 s 6882 40227 6980 40325 4 vdd
rlabel metal3 s 6882 33549 6980 33647 4 vdd
rlabel metal3 s 7660 741 7758 839 4 vdd
rlabel metal3 s 6882 3887 6980 3985 4 vdd
rlabel metal3 s 6450 19687 6548 19785 4 vdd
rlabel metal3 s 7660 26416 7758 26514 4 vdd
rlabel metal3 s 6882 10639 6980 10737 4 vdd
rlabel metal3 s 6450 2739 6548 2837 4 vdd
rlabel metal3 s 7660 4691 7758 4789 4 vdd
rlabel metal3 s 6450 33117 6548 33215 4 vdd
rlabel metal3 s 7660 39846 7758 39944 4 vdd
rlabel metal3 s 6450 13009 6548 13107 4 vdd
rlabel metal3 s 6882 24069 6980 24167 4 vdd
rlabel metal3 s 7660 30761 7758 30859 4 vdd
rlabel metal3 s 6882 44609 6980 44707 4 vdd
rlabel metal3 s 6882 41017 6980 41115 4 vdd
rlabel metal3 s 6450 33907 6548 34005 4 vdd
rlabel metal3 s 7660 6271 7758 6369 4 vdd
rlabel metal3 s 6450 43387 6548 43485 4 vdd
rlabel metal3 s 7660 18911 7758 19009 4 vdd
rlabel metal3 s 6882 38289 6980 38387 4 vdd
rlabel metal3 s 6450 4677 6548 4775 4 vdd
rlabel metal3 s 7660 4296 7758 4394 4 vdd
rlabel metal3 s 6450 17749 6548 17847 4 vdd
rlabel metal3 s 7660 3111 7758 3209 4 vdd
rlabel metal3 s 6450 20477 6548 20575 4 vdd
rlabel metal3 s 6882 4319 6980 4417 4 vdd
rlabel metal3 s 7660 29971 7758 30069 4 vdd
rlabel metal3 s 7660 5876 7758 5974 4 vdd
rlabel metal3 s 6450 35487 6548 35585 4 vdd
rlabel metal3 s 7660 46166 7758 46264 4 vdd
rlabel metal3 s 6882 16527 6980 16625 4 vdd
rlabel metal3 s 6882 42597 6980 42695 4 vdd
rlabel metal3 s 6450 11429 6548 11527 4 vdd
rlabel metal3 s 7660 43006 7758 43104 4 vdd
rlabel metal3 s 6450 23279 6548 23377 4 vdd
rlabel metal3 s 6882 40659 6980 40757 4 vdd
rlabel metal3 s 6882 3529 6980 3627 4 vdd
rlabel metal3 s 6450 22847 6548 22945 4 vdd
rlabel metal3 s 3468 5899 3566 5997 4 vdd
rlabel metal3 s 6882 11429 6980 11527 4 vdd
rlabel metal3 s 6450 43029 6548 43127 4 vdd
rlabel metal3 s 3036 7479 3134 7577 4 vdd
rlabel metal3 s 7660 29576 7758 29674 4 vdd
rlabel metal3 s 7660 49326 7758 49424 4 vdd
rlabel metal3 s 7660 14961 7758 15059 4 vdd
rlabel metal3 s 6882 48127 6980 48225 4 vdd
rlabel metal3 s 6450 48917 6548 49015 4 vdd
rlabel metal3 s 6450 32327 6548 32425 4 vdd
rlabel metal3 s 6450 3097 6548 3195 4 vdd
rlabel metal3 s 6882 20477 6980 20575 4 vdd
rlabel metal3 s 6450 35919 6548 36017 4 vdd
rlabel metal3 s 6882 44967 6980 45065 4 vdd
rlabel metal3 s 6450 6257 6548 6355 4 vdd
rlabel metal3 s 6882 19687 6980 19785 4 vdd
rlabel metal3 s 6450 7479 6548 7577 4 vdd
rlabel metal3 s 6882 10207 6980 10305 4 vdd
rlabel metal3 s 6882 31969 6980 32067 4 vdd
rlabel metal3 s 6882 1517 6980 1615 4 vdd
rlabel metal3 s 6450 38647 6548 38745 4 vdd
rlabel metal3 s 6450 44609 6548 44707 4 vdd
rlabel metal3 s 6450 42239 6548 42337 4 vdd
rlabel metal3 s 4246 3506 4344 3604 4 vdd
rlabel metal3 s 6450 12219 6548 12317 4 vdd
rlabel metal3 s 6882 28377 6980 28475 4 vdd
rlabel metal3 s 6450 20909 6548 21007 4 vdd
rlabel metal3 s 6450 47337 6548 47435 4 vdd
rlabel metal3 s 7660 45376 7758 45474 4 vdd
rlabel metal3 s 7660 44586 7758 44684 4 vdd
rlabel metal3 s 7660 38661 7758 38759 4 vdd
rlabel metal3 s 6450 9849 6548 9947 4 vdd
rlabel metal3 s 6882 8627 6980 8725 4 vdd
rlabel metal3 s 7660 16541 7758 16639 4 vdd
rlabel metal3 s 6882 30747 6980 30845 4 vdd
rlabel metal3 s 6450 14947 6548 15045 4 vdd
rlabel metal3 s 7660 50116 7758 50214 4 vdd
rlabel metal3 s 6882 22057 6980 22155 4 vdd
rlabel metal3 s 6882 9417 6980 9515 4 vdd
rlabel metal3 s 6450 49349 6548 49447 4 vdd
rlabel metal3 s 6450 15379 6548 15477 4 vdd
rlabel metal3 s 6450 10639 6548 10737 4 vdd
rlabel metal3 s 7660 37476 7758 37574 4 vdd
rlabel metal3 s 6450 35129 6548 35227 4 vdd
rlabel metal3 s 6450 20119 6548 20217 4 vdd
rlabel metal3 s 6450 26797 6548 26895 4 vdd
rlabel metal3 s 7660 22466 7758 22564 4 vdd
rlabel metal3 s 6450 34697 6548 34795 4 vdd
rlabel metal3 s 6450 44967 6548 45065 4 vdd
rlabel metal3 s 7660 35106 7758 35204 4 vdd
rlabel metal3 s 7660 41426 7758 41524 4 vdd
rlabel metal3 s 6882 31537 6980 31635 4 vdd
rlabel metal3 s 6882 27229 6980 27327 4 vdd
rlabel metal3 s 7660 10616 7758 10714 4 vdd
rlabel metal3 s 6882 33117 6980 33215 4 vdd
rlabel metal3 s 6450 18897 6548 18995 4 vdd
rlabel metal3 s 7660 35501 7758 35599 4 vdd
rlabel metal3 s 6882 16959 6980 17057 4 vdd
rlabel metal3 s 2148 346 2246 444 4 vdd
rlabel metal3 s 7660 37081 7758 37179 4 vdd
rlabel metal3 s 6882 13009 6980 13107 4 vdd
rlabel metal3 s 6882 35919 6980 36017 4 vdd
rlabel metal3 s 6882 8269 6980 8367 4 vdd
rlabel metal3 s 6450 7837 6548 7935 4 vdd
rlabel metal3 s 7660 43796 7758 43894 4 vdd
rlabel metal3 s 7660 8641 7758 8739 4 vdd
rlabel metal3 s 4246 7456 4344 7554 4 vdd
rlabel metal3 s 3468 6689 3566 6787 4 vdd
rlabel metal3 s 6450 8627 6548 8725 4 vdd
rlabel metal3 s 6450 26439 6548 26537 4 vdd
rlabel metal3 s 6882 10997 6980 11095 4 vdd
rlabel metal3 s 6882 20909 6980 21007 4 vdd
rlabel metal3 s 7660 11406 7758 11504 4 vdd
rlabel metal3 s 6882 3097 6980 3195 4 vdd
rlabel metal3 s 6450 25649 6548 25747 4 vdd
rlabel metal3 s 6882 39079 6980 39177 4 vdd
rlabel metal3 s 7660 18516 7758 18614 4 vdd
rlabel metal3 s 6882 6689 6980 6787 4 vdd
rlabel metal3 s 3468 5109 3566 5207 4 vdd
rlabel metal3 s 3471 2723 3569 2821 4 vdd
rlabel metal3 s 6450 18539 6548 18637 4 vdd
rlabel metal3 s 6882 32759 6980 32857 4 vdd
rlabel metal3 s 7660 15356 7758 15454 4 vdd
rlabel metal3 s 6882 46979 6980 47077 4 vdd
rlabel metal3 s 6450 36709 6548 36807 4 vdd
rlabel metal3 s 7660 21281 7758 21379 4 vdd
rlabel metal3 s 7660 36686 7758 36784 4 vdd
rlabel metal3 s 6450 30389 6548 30487 4 vdd
rlabel metal3 s 6450 27587 6548 27685 4 vdd
rlabel metal3 s 6882 13367 6980 13465 4 vdd
rlabel metal3 s 6450 27229 6548 27327 4 vdd
rlabel metal3 s 4246 1136 4344 1234 4 vdd
rlabel metal3 s 6450 39437 6548 39535 4 vdd
rlabel metal3 s 6450 14589 6548 14687 4 vdd
rlabel metal3 s 7660 18121 7758 18219 4 vdd
rlabel metal3 s 6450 16169 6548 16267 4 vdd
rlabel metal3 s 7660 9431 7758 9529 4 vdd
rlabel metal3 s 7660 20886 7758 20984 4 vdd
rlabel metal3 s 6450 3887 6548 3985 4 vdd
rlabel metal3 s 7660 48536 7758 48634 4 vdd
rlabel metal3 s 6882 13799 6980 13897 4 vdd
rlabel metal3 s 6450 31179 6548 31277 4 vdd
rlabel metal3 s 7660 7851 7758 7949 4 vdd
rlabel metal3 s 7660 12196 7758 12294 4 vdd
rlabel metal3 s 7660 37871 7758 37969 4 vdd
rlabel metal3 s 6882 23637 6980 23735 4 vdd
rlabel metal3 s 7660 44191 7758 44289 4 vdd
rlabel metal3 s 6882 36277 6980 36375 4 vdd
rlabel metal3 s 7660 9036 7758 9134 4 vdd
rlabel metal3 s 7660 49721 7758 49819 4 vdd
rlabel metal3 s 7660 5481 7758 5579 4 vdd
rlabel metal3 s 6882 12219 6980 12317 4 vdd
rlabel metal3 s 6882 29167 6980 29265 4 vdd
rlabel metal3 s 6450 10997 6548 11095 4 vdd
rlabel metal3 s 3036 5109 3134 5207 4 vdd
rlabel metal3 s 7660 29181 7758 29279 4 vdd
rlabel metal3 s 7660 10221 7758 10319 4 vdd
rlabel metal3 s 7660 41821 7758 41919 4 vdd
rlabel metal3 s 6882 369 6980 467 4 vdd
rlabel metal3 s 6882 7047 6980 7145 4 vdd
rlabel metal3 s 6882 44177 6980 44275 4 vdd
rlabel metal3 s 6882 47769 6980 47867 4 vdd
rlabel metal3 s 6450 21267 6548 21365 4 vdd
rlabel metal3 s 6882 14589 6980 14687 4 vdd
rlabel metal3 s 6882 42239 6980 42337 4 vdd
rlabel metal3 s 7660 22071 7758 22169 4 vdd
rlabel metal3 s 7660 38266 7758 38364 4 vdd
rlabel metal3 s 7660 2716 7758 2814 4 vdd
rlabel metal3 s 6450 34339 6548 34437 4 vdd
rlabel metal3 s 6450 48559 6548 48657 4 vdd
rlabel metal3 s 7660 19701 7758 19799 4 vdd
rlabel metal3 s 7660 26021 7758 26119 4 vdd
rlabel metal3 s 6450 40659 6548 40757 4 vdd
rlabel metal3 s 6882 727 6980 825 4 vdd
rlabel metal3 s 3468 7479 3566 7577 4 vdd
rlabel metal3 s 7660 14566 7758 14664 4 vdd
rlabel metal3 s 6882 25217 6980 25315 4 vdd
rlabel metal3 s 6450 28019 6548 28117 4 vdd
rlabel metal3 s 6450 3529 6548 3627 4 vdd
rlabel metal3 s 6450 47769 6548 47867 4 vdd
rlabel metal3 s 6882 29599 6980 29697 4 vdd
rlabel metal3 s 6882 30389 6980 30487 4 vdd
rlabel metal3 s 6450 31969 6548 32067 4 vdd
rlabel metal3 s 6882 39869 6980 39967 4 vdd
port 136 se
rlabel metal3 s 7264 35501 7362 35599 4 gnd
rlabel metal3 s 6025 41449 6123 41547 4 gnd
rlabel metal3 s 7264 19306 7362 19404 4 gnd
rlabel metal3 s 3046 2723 3144 2821 4 gnd
rlabel metal3 s 7264 14171 7362 14269 4 gnd
rlabel metal3 s 6025 21325 6123 21423 4 gnd
rlabel metal3 s 6025 48185 6123 48283 4 gnd
rlabel metal3 s 6025 7105 6123 7203 4 gnd
rlabel metal3 s 7264 21676 7362 21774 4 gnd
rlabel metal3 s 7264 36291 7362 36389 4 gnd
rlabel metal3 s 6025 30015 6123 30113 4 gnd
rlabel metal3 s 6025 43029 6123 43127 4 gnd
rlabel metal3 s 7264 12591 7362 12689 4 gnd
rlabel metal3 s 7264 43006 7362 43104 4 gnd
rlabel metal3 s 6025 18539 6123 18637 4 gnd
rlabel metal3 s 7264 26416 7362 26514 4 gnd
rlabel metal3 s 7264 3506 7362 3604 4 gnd
rlabel metal3 s 6025 24859 6123 24957 4 gnd
rlabel metal3 s 6025 39079 6123 39177 4 gnd
rlabel metal3 s 6025 2365 6123 2463 4 gnd
rlabel metal3 s 6025 23279 6123 23377 4 gnd
rlabel metal3 s 6025 34755 6123 34853 4 gnd
rlabel metal3 s 6025 43819 6123 43917 4 gnd
rlabel metal3 s 6025 50139 6123 50237 4 gnd
rlabel metal3 s 7264 48536 7362 48634 4 gnd
rlabel metal3 s 6025 10265 6123 10363 4 gnd
rlabel metal3 s 6025 11055 6123 11153 4 gnd
rlabel metal3 s 7264 18516 7362 18614 4 gnd
rlabel metal3 s 7264 39056 7362 39154 4 gnd
rlabel metal3 s 7264 30366 7362 30464 4 gnd
rlabel metal3 s 6025 46189 6123 46287 4 gnd
rlabel metal3 s 6025 48975 6123 49073 4 gnd
rlabel metal3 s 7264 32341 7362 32439 4 gnd
rlabel metal3 s 6025 17375 6123 17473 4 gnd
rlabel metal3 s 6025 20909 6123 21007 4 gnd
rlabel metal3 s 7264 10221 7362 10319 4 gnd
rlabel metal3 s 7264 33921 7362 34019 4 gnd
rlabel metal3 s 7264 39451 7362 39549 4 gnd
rlabel metal3 s 7264 25231 7362 25329 4 gnd
rlabel metal3 s 7264 42216 7362 42314 4 gnd
rlabel metal3 s 6025 29225 6123 29323 4 gnd
rlabel metal3 s 6025 32385 6123 32483 4 gnd
rlabel metal3 s 7264 46166 7362 46264 4 gnd
rlabel metal3 s 7264 20491 7362 20589 4 gnd
rlabel metal3 s 6025 42655 6123 42753 4 gnd
rlabel metal3 s 6025 24069 6123 24167 4 gnd
rlabel metal3 s 6025 48559 6123 48657 4 gnd
rlabel metal3 s 6025 49349 6123 49447 4 gnd
rlabel metal3 s 6025 785 6123 883 4 gnd
rlabel metal3 s 6025 21699 6123 21797 4 gnd
rlabel metal3 s 7264 34316 7362 34414 4 gnd
rlabel metal3 s 6025 29599 6123 29697 4 gnd
rlabel metal3 s 7264 16541 7362 16639 4 gnd
rlabel metal3 s 3046 353 3144 451 4 gnd
rlabel metal3 s 2611 5109 2709 5207 4 gnd
rlabel metal3 s 6025 20535 6123 20633 4 gnd
rlabel metal3 s 7264 8246 7362 8344 4 gnd
rlabel metal3 s 6025 42239 6123 42337 4 gnd
rlabel metal3 s 2611 7479 2709 7577 4 gnd
rlabel metal3 s 6025 9059 6123 9157 4 gnd
rlabel metal3 s 7264 38661 7362 38759 4 gnd
rlabel metal3 s 6025 32759 6123 32857 4 gnd
rlabel metal3 s 7264 26811 7362 26909 4 gnd
rlabel metal3 s 7264 44981 7362 45079 4 gnd
rlabel metal3 s 6025 30805 6123 30903 4 gnd
rlabel metal3 s 7264 741 7362 839 4 gnd
rlabel metal3 s 6025 3529 6123 3627 4 gnd
rlabel metal3 s 3850 1136 3948 1234 4 gnd
rlabel metal3 s 2611 5899 2709 5997 4 gnd
rlabel metal3 s 6025 8269 6123 8367 4 gnd
rlabel metal3 s 7264 48141 7362 48239 4 gnd
rlabel metal3 s 7264 36686 7362 36784 4 gnd
rlabel metal3 s 7264 7456 7362 7554 4 gnd
rlabel metal3 s 3850 5086 3948 5184 4 gnd
rlabel metal3 s 6025 28435 6123 28533 4 gnd
rlabel metal3 s 7264 41821 7362 41919 4 gnd
rlabel metal3 s 7264 45376 7362 45474 4 gnd
rlabel metal3 s 6025 36335 6123 36433 4 gnd
rlabel metal3 s 7264 6271 7362 6369 4 gnd
rlabel metal3 s 7264 15356 7362 15454 4 gnd
rlabel metal3 s 7264 3901 7362 3999 4 gnd
rlabel metal3 s 6025 18955 6123 19053 4 gnd
rlabel metal3 s 7264 1136 7362 1234 4 gnd
rlabel metal3 s 7264 14566 7362 14664 4 gnd
rlabel metal3 s 7264 24441 7362 24539 4 gnd
rlabel metal3 s 7264 16146 7362 16244 4 gnd
rlabel metal3 s 6025 23695 6123 23793 4 gnd
rlabel metal3 s 7264 12196 7362 12294 4 gnd
rlabel metal3 s 2611 6689 2709 6787 4 gnd
rlabel metal3 s 6025 37915 6123 38013 4 gnd
rlabel metal3 s 6025 20119 6123 20217 4 gnd
rlabel metal3 s 7264 8641 7362 8739 4 gnd
rlabel metal3 s 7264 9826 7362 9924 4 gnd
rlabel metal3 s 7264 20096 7362 20194 4 gnd
rlabel metal3 s 6025 28809 6123 28907 4 gnd
rlabel metal3 s 6025 47395 6123 47493 4 gnd
rlabel metal3 s 6025 27645 6123 27743 4 gnd
rlabel metal3 s 6025 39869 6123 39967 4 gnd
rlabel metal3 s 7264 17331 7362 17429 4 gnd
rlabel metal3 s 6025 15795 6123 15893 4 gnd
rlabel metal3 s 7264 37081 7362 37179 4 gnd
rlabel metal3 s 7264 35896 7362 35994 4 gnd
rlabel metal3 s 6025 26065 6123 26163 4 gnd
rlabel metal3 s 6025 13425 6123 13523 4 gnd
rlabel metal3 s 7264 13776 7362 13874 4 gnd
rlabel metal3 s 6025 43445 6123 43543 4 gnd
rlabel metal3 s 7264 18121 7362 18219 4 gnd
rlabel metal3 s 7264 5086 7362 5184 4 gnd
rlabel metal3 s 7264 15751 7362 15849 4 gnd
rlabel metal3 s 7264 22071 7362 22169 4 gnd
rlabel metal3 s 6025 31969 6123 32067 4 gnd
rlabel metal3 s 7264 22861 7362 22959 4 gnd
rlabel metal3 s 6025 12219 6123 12317 4 gnd
rlabel metal3 s 6025 11429 6123 11527 4 gnd
rlabel metal3 s 6025 2739 6123 2837 4 gnd
rlabel metal3 s 6025 16169 6123 16267 4 gnd
rlabel metal3 s 6025 37499 6123 37597 4 gnd
rlabel metal3 s 6025 41075 6123 41173 4 gnd
rlabel metal3 s 6025 9475 6123 9573 4 gnd
rlabel metal3 s 7264 43796 7362 43894 4 gnd
rlabel metal3 s 6025 9849 6123 9947 4 gnd
rlabel metal3 s 3850 7456 3948 7554 4 gnd
rlabel metal3 s 7264 3111 7362 3209 4 gnd
rlabel metal3 s 6025 35129 6123 35227 4 gnd
rlabel metal3 s 6025 47769 6123 47867 4 gnd
rlabel metal3 s 6025 49765 6123 49863 4 gnd
rlabel metal3 s 7264 11406 7362 11504 4 gnd
rlabel metal3 s 6025 13009 6123 13107 4 gnd
rlabel metal3 s 6025 26855 6123 26953 4 gnd
rlabel metal3 s 7264 45771 7362 45869 4 gnd
rlabel metal3 s 6025 1159 6123 1257 4 gnd
rlabel metal3 s 6025 13799 6123 13897 4 gnd
rlabel metal3 s 6025 15379 6123 15477 4 gnd
rlabel metal3 s 6025 1575 6123 1673 4 gnd
rlabel metal3 s 7264 24046 7362 24144 4 gnd
rlabel metal3 s 6025 39495 6123 39593 4 gnd
rlabel metal3 s 6025 12635 6123 12733 4 gnd
rlabel metal3 s 7264 12986 7362 13084 4 gnd
rlabel metal3 s 3850 346 3948 444 4 gnd
rlabel metal3 s 6025 38705 6123 38803 4 gnd
rlabel metal3 s 6025 46605 6123 46703 4 gnd
rlabel metal3 s 6025 31179 6123 31277 4 gnd
rlabel metal3 s 7264 30761 7362 30859 4 gnd
rlabel metal3 s 7264 13381 7362 13479 4 gnd
rlabel metal3 s 6025 5109 6123 5207 4 gnd
rlabel metal3 s 7264 44586 7362 44684 4 gnd
rlabel metal3 s 6025 24485 6123 24583 4 gnd
rlabel metal3 s 3850 2716 3948 2814 4 gnd
rlabel metal3 s 7264 20886 7362 20984 4 gnd
rlabel metal3 s 6025 7895 6123 7993 4 gnd
rlabel metal3 s 6025 17749 6123 17847 4 gnd
rlabel metal3 s 7264 27601 7362 27699 4 gnd
rlabel metal3 s 7264 38266 7362 38364 4 gnd
rlabel metal3 s 6025 22115 6123 22213 4 gnd
rlabel metal3 s 6025 30389 6123 30487 4 gnd
rlabel metal3 s 3850 5876 3948 5974 4 gnd
rlabel metal3 s 6025 25649 6123 25747 4 gnd
rlabel metal3 s 7264 25626 7362 25724 4 gnd
rlabel metal3 s 7264 16936 7362 17034 4 gnd
rlabel metal3 s 7264 42611 7362 42709 4 gnd
rlabel metal3 s 6025 36709 6123 36807 4 gnd
rlabel metal3 s 7264 43401 7362 43499 4 gnd
rlabel metal3 s 6025 16585 6123 16683 4 gnd
rlabel metal3 s 7264 29576 7362 29674 4 gnd
rlabel metal3 s 6025 34339 6123 34437 4 gnd
rlabel metal3 s 6025 44235 6123 44333 4 gnd
rlabel metal3 s 1752 346 1850 444 4 gnd
rlabel metal3 s 7264 7851 7362 7949 4 gnd
rlabel metal3 s 7264 29181 7362 29279 4 gnd
rlabel metal3 s 6025 25275 6123 25373 4 gnd
rlabel metal3 s 6025 33549 6123 33647 4 gnd
rlabel metal3 s 7264 48931 7362 49029 4 gnd
rlabel metal3 s 6025 46979 6123 47077 4 gnd
rlabel metal3 s 7264 11011 7362 11109 4 gnd
rlabel metal3 s 7264 23256 7362 23354 4 gnd
rlabel metal3 s 7264 22466 7362 22564 4 gnd
rlabel metal3 s 6025 45815 6123 45913 4 gnd
rlabel metal3 s 7264 26021 7362 26119 4 gnd
rlabel metal3 s 1156 5086 1254 5184 4 gnd
rlabel metal3 s 7264 2716 7362 2814 4 gnd
rlabel metal3 s 6025 3155 6123 3253 4 gnd
rlabel metal3 s 7264 41426 7362 41524 4 gnd
rlabel metal3 s 7264 346 7362 444 4 gnd
rlabel metal3 s 3850 6666 3948 6764 4 gnd
rlabel metal3 s 7264 31946 7362 32044 4 gnd
rlabel metal3 s 6025 37125 6123 37223 4 gnd
rlabel metal3 s 7264 27206 7362 27304 4 gnd
rlabel metal3 s 6025 1949 6123 2047 4 gnd
rlabel metal3 s 6025 6689 6123 6787 4 gnd
rlabel metal3 s 7264 40636 7362 40734 4 gnd
rlabel metal3 s 7264 46956 7362 47054 4 gnd
rlabel metal3 s 7264 6666 7362 6764 4 gnd
rlabel metal3 s 7264 18911 7362 19009 4 gnd
rlabel metal3 s 6025 16959 6123 17057 4 gnd
rlabel metal3 s 7264 32736 7362 32834 4 gnd
rlabel metal3 s 7264 1926 7362 2024 4 gnd
rlabel metal3 s 7264 7061 7362 7159 4 gnd
rlabel metal3 s 7264 10616 7362 10714 4 gnd
rlabel metal3 s 6025 369 6123 467 4 gnd
rlabel metal3 s 7264 11801 7362 11899 4 gnd
rlabel metal3 s 7264 28391 7362 28489 4 gnd
rlabel metal3 s 7264 49721 7362 49819 4 gnd
rlabel metal3 s 7264 17726 7362 17824 4 gnd
rlabel metal3 s 7264 33526 7362 33624 4 gnd
rlabel metal3 s 6025 41865 6123 41963 4 gnd
rlabel metal3 s 7264 41031 7362 41129 4 gnd
rlabel metal3 s 6025 22489 6123 22587 4 gnd
rlabel metal3 s 6025 40659 6123 40757 4 gnd
rlabel metal3 s 7264 47746 7362 47844 4 gnd
rlabel metal3 s 6025 7479 6123 7577 4 gnd
rlabel metal3 s 3046 3513 3144 3611 4 gnd
rlabel metal3 s 7264 34711 7362 34809 4 gnd
rlabel metal3 s 6025 19745 6123 19843 4 gnd
rlabel metal3 s 6025 35545 6123 35643 4 gnd
rlabel metal3 s 7264 28786 7362 28884 4 gnd
rlabel metal3 s 7264 31551 7362 31649 4 gnd
rlabel metal3 s 7264 39846 7362 39944 4 gnd
rlabel metal3 s 7264 47351 7362 47449 4 gnd
rlabel metal3 s 7264 40241 7362 40339 4 gnd
rlabel metal3 s 7264 31156 7362 31254 4 gnd
rlabel metal3 s 7264 14961 7362 15059 4 gnd
rlabel metal3 s 1752 2716 1850 2814 4 gnd
rlabel metal3 s 7264 5876 7362 5974 4 gnd
rlabel metal3 s 6025 4319 6123 4417 4 gnd
rlabel metal3 s 6025 15005 6123 15103 4 gnd
rlabel metal3 s 6025 26439 6123 26537 4 gnd
rlabel metal3 s 7264 37871 7362 37969 4 gnd
rlabel metal3 s 6025 35919 6123 36017 4 gnd
rlabel metal3 s 6025 5899 6123 5997 4 gnd
rlabel metal3 s 7264 2321 7362 2419 4 gnd
rlabel metal3 s 7264 50116 7362 50214 4 gnd
rlabel metal3 s 7264 33131 7362 33229 4 gnd
rlabel metal3 s 6025 22905 6123 23003 4 gnd
rlabel metal3 s 6025 38289 6123 38387 4 gnd
rlabel metal3 s 6025 40285 6123 40383 4 gnd
rlabel metal3 s 6025 14215 6123 14313 4 gnd
rlabel metal3 s 7264 19701 7362 19799 4 gnd
rlabel metal3 s 7264 4296 7362 4394 4 gnd
rlabel metal3 s 7264 29971 7362 30069 4 gnd
rlabel metal3 s 6025 45025 6123 45123 4 gnd
rlabel metal3 s 7264 49326 7362 49424 4 gnd
rlabel metal3 s 6025 11845 6123 11943 4 gnd
rlabel metal3 s 6025 33965 6123 34063 4 gnd
rlabel metal3 s 7264 9431 7362 9529 4 gnd
rlabel metal3 s 6025 45399 6123 45497 4 gnd
rlabel metal3 s 7264 37476 7362 37574 4 gnd
rlabel metal3 s 6025 8685 6123 8783 4 gnd
rlabel metal3 s 6025 27229 6123 27327 4 gnd
rlabel metal3 s 7264 44191 7362 44289 4 gnd
rlabel metal3 s 7264 35106 7362 35204 4 gnd
rlabel metal3 s 7264 46561 7362 46659 4 gnd
rlabel metal3 s 6025 4735 6123 4833 4 gnd
rlabel metal3 s 6025 28019 6123 28117 4 gnd
rlabel metal3 s 6025 5525 6123 5623 4 gnd
rlabel metal3 s 6025 6315 6123 6413 4 gnd
rlabel metal3 s 7264 21281 7362 21379 4 gnd
rlabel metal3 s 6025 33175 6123 33273 4 gnd
rlabel metal3 s 6025 19329 6123 19427 4 gnd
rlabel metal3 s 6025 44609 6123 44707 4 gnd
rlabel metal3 s 7264 24836 7362 24934 4 gnd
rlabel metal3 s 6025 10639 6123 10737 4 gnd
rlabel metal3 s 7264 5481 7362 5579 4 gnd
rlabel metal3 s 7264 23651 7362 23749 4 gnd
rlabel metal3 s 7264 1531 7362 1629 4 gnd
rlabel metal3 s 6025 31595 6123 31693 4 gnd
rlabel metal3 s 7264 4691 7362 4789 4 gnd
rlabel metal3 s 3046 1143 3144 1241 4 gnd
rlabel metal3 s 6025 18165 6123 18263 4 gnd
rlabel metal3 s 7264 27996 7362 28094 4 gnd
rlabel metal3 s 3850 3506 3948 3604 4 gnd
rlabel metal3 s 6025 3945 6123 4043 4 gnd
rlabel metal3 s 6025 14589 6123 14687 4 gnd
rlabel metal3 s 7264 9036 7362 9134 4 gnd
port 137 se
<< properties >>
string FIXED_BBOX 4505 -32 4569 0
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 8759706
string GDS_START 8451404
<< end >>
