magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1443 -1243 1078 1278
<< labels >>
flabel comment s -183 17 -183 17 0 FreeSans 1000 0 0 0 LI_JUMPER_OK
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36328718
string GDS_START 36326450
<< end >>
