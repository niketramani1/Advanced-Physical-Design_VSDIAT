magic
tech sky130A
magscale 1 2
timestamp 1624855595
<< checkpaint >>
rect -1298 -1308 2678 1852
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 543 47 573 119
rect 629 47 659 119
rect 724 47 754 131
rect 921 47 951 177
rect 1008 47 1038 177
rect 1092 47 1122 177
rect 1183 47 1213 177
rect 1271 47 1301 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 652 413 682 497
rect 724 413 754 497
rect 921 297 951 497
rect 1008 297 1038 497
rect 1092 297 1122 497
rect 1183 297 1213 497
rect 1271 297 1301 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 869 133 921 177
rect 674 119 724 131
rect 465 47 543 119
rect 573 107 629 119
rect 573 73 584 107
rect 618 73 629 107
rect 573 47 629 73
rect 659 47 724 119
rect 754 106 806 131
rect 754 72 764 106
rect 798 72 806 106
rect 754 47 806 72
rect 869 99 877 133
rect 911 99 921 133
rect 869 47 921 99
rect 951 127 1008 177
rect 951 93 964 127
rect 998 93 1008 127
rect 951 47 1008 93
rect 1038 133 1092 177
rect 1038 99 1048 133
rect 1082 99 1092 133
rect 1038 47 1092 99
rect 1122 127 1183 177
rect 1122 93 1139 127
rect 1173 93 1183 127
rect 1122 47 1183 93
rect 1213 127 1271 177
rect 1213 93 1223 127
rect 1257 93 1271 127
rect 1213 47 1271 93
rect 1301 127 1353 177
rect 1301 93 1311 127
rect 1345 93 1353 127
rect 1301 47 1353 93
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 652 497
rect 561 451 596 485
rect 630 451 652 485
rect 561 413 652 451
rect 682 413 724 497
rect 754 477 806 497
rect 754 443 764 477
rect 798 443 806 477
rect 754 413 806 443
rect 869 471 921 497
rect 869 437 877 471
rect 911 437 921 471
rect 465 369 515 413
rect 869 368 921 437
rect 869 334 877 368
rect 911 334 921 368
rect 869 297 921 334
rect 951 484 1008 497
rect 951 450 964 484
rect 998 450 1008 484
rect 951 364 1008 450
rect 951 330 964 364
rect 998 330 1008 364
rect 951 297 1008 330
rect 1038 475 1092 497
rect 1038 441 1048 475
rect 1082 441 1092 475
rect 1038 384 1092 441
rect 1038 350 1048 384
rect 1082 350 1092 384
rect 1038 297 1092 350
rect 1122 475 1183 497
rect 1122 441 1139 475
rect 1173 441 1183 475
rect 1122 384 1183 441
rect 1122 350 1139 384
rect 1173 350 1183 384
rect 1122 297 1183 350
rect 1213 475 1271 497
rect 1213 441 1223 475
rect 1257 441 1271 475
rect 1213 384 1271 441
rect 1213 350 1223 384
rect 1257 350 1271 384
rect 1213 297 1271 350
rect 1301 475 1353 497
rect 1301 441 1311 475
rect 1345 441 1353 475
rect 1301 384 1353 441
rect 1301 350 1311 384
rect 1345 350 1353 384
rect 1301 297 1353 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 584 73 618 107
rect 764 72 798 106
rect 877 99 911 133
rect 964 93 998 127
rect 1048 99 1082 133
rect 1139 93 1173 127
rect 1223 93 1257 127
rect 1311 93 1345 127
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 596 451 630 485
rect 764 443 798 477
rect 877 437 911 471
rect 877 334 911 368
rect 964 450 998 484
rect 964 330 998 364
rect 1048 441 1082 475
rect 1048 350 1082 384
rect 1139 441 1173 475
rect 1139 350 1173 384
rect 1223 441 1257 475
rect 1223 350 1257 384
rect 1311 441 1345 475
rect 1311 350 1345 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 652 497 682 523
rect 724 497 754 523
rect 921 497 951 523
rect 1008 497 1038 523
rect 1092 497 1122 523
rect 1183 497 1213 523
rect 1271 497 1301 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 652 375 682 413
rect 507 321 561 337
rect 603 365 682 375
rect 603 331 619 365
rect 653 331 682 365
rect 603 321 682 331
rect 724 373 754 413
rect 724 357 812 373
rect 724 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 507 279 561 287
rect 724 307 812 323
rect 507 271 659 279
rect 531 249 659 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 533 191 587 207
rect 533 157 543 191
rect 577 157 587 191
rect 435 131 465 153
rect 533 141 587 157
rect 543 119 573 141
rect 629 119 659 249
rect 724 131 754 307
rect 921 265 951 297
rect 1008 265 1038 297
rect 1092 265 1122 297
rect 1183 265 1213 297
rect 1271 265 1301 297
rect 796 249 951 265
rect 796 215 806 249
rect 840 215 951 249
rect 796 199 951 215
rect 993 249 1301 265
rect 993 215 1003 249
rect 1037 215 1301 249
rect 993 199 1301 215
rect 921 177 951 199
rect 1008 177 1038 199
rect 1092 177 1122 199
rect 1183 177 1213 199
rect 1271 177 1301 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 543 21 573 47
rect 629 21 659 47
rect 724 21 754 47
rect 921 21 951 47
rect 1008 21 1038 47
rect 1092 21 1122 47
rect 1183 21 1213 47
rect 1271 21 1301 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 543 157 577 191
rect 806 215 840 249
rect 1003 215 1037 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 580 451 596 485
rect 630 451 730 485
rect 391 417 454 451
rect 425 383 454 417
rect 391 367 454 383
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 321 551 357
rect 494 287 517 321
rect 494 271 551 287
rect 585 365 653 399
rect 585 331 619 365
rect 585 323 653 331
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 394 203 468 219
rect 585 207 619 283
rect 696 265 730 451
rect 764 477 824 527
rect 798 443 824 477
rect 764 427 824 443
rect 877 471 921 487
rect 911 437 921 471
rect 877 373 921 437
rect 768 368 921 373
rect 768 357 877 368
rect 802 334 877 357
rect 911 334 921 368
rect 802 323 921 334
rect 768 307 921 323
rect 887 265 921 307
rect 957 484 1014 527
rect 957 450 964 484
rect 998 450 1014 484
rect 957 364 1014 450
rect 957 330 964 364
rect 998 330 1014 364
rect 957 299 1014 330
rect 1048 475 1105 491
rect 1082 441 1105 475
rect 1048 384 1105 441
rect 1082 350 1105 384
rect 1048 299 1105 350
rect 1139 475 1189 527
rect 1173 441 1189 475
rect 1139 384 1189 441
rect 1173 350 1189 384
rect 1139 299 1189 350
rect 1223 475 1277 491
rect 1257 441 1277 475
rect 1223 384 1277 441
rect 1257 350 1277 384
rect 1071 265 1105 299
rect 1223 265 1277 350
rect 1311 475 1363 527
rect 1345 441 1363 475
rect 1311 384 1363 441
rect 1345 350 1363 384
rect 1311 299 1363 350
rect 696 249 840 265
rect 696 233 806 249
rect 394 169 434 203
rect 394 157 468 169
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 543 191 619 207
rect 577 157 619 191
rect 307 123 428 153
rect 543 141 619 157
rect 666 215 806 233
rect 666 199 840 215
rect 887 249 1037 265
rect 887 215 1003 249
rect 887 199 1037 215
rect 1071 199 1363 265
rect 307 119 341 123
rect 666 107 700 199
rect 887 149 921 199
rect 1071 149 1105 199
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 568 73 584 107
rect 618 73 700 107
rect 877 133 921 149
rect 375 17 441 55
rect 748 72 764 106
rect 798 72 814 106
rect 911 99 921 133
rect 877 83 921 99
rect 957 127 1014 143
rect 957 93 964 127
rect 998 93 1014 127
rect 748 17 814 72
rect 957 17 1014 93
rect 1048 133 1105 149
rect 1082 99 1105 133
rect 1048 83 1105 99
rect 1139 127 1189 165
rect 1173 93 1189 127
rect 1139 17 1189 93
rect 1223 127 1277 199
rect 1257 93 1277 127
rect 1223 77 1277 93
rect 1311 127 1363 143
rect 1345 93 1363 127
rect 1311 17 1363 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 494 357 528 391
rect 586 289 620 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1059 357 1093 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1059 425 1093 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1059 85 1093 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1140 221 1174 255 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1232 221 1266 255 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1324 221 1358 255 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1243 357 1277 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1243 425 1277 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1243 153 1277 187 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1243 85 1277 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 dlxtn_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2381050
string GDS_START 2369358
string path 0.000 13.600 34.500 13.600 
<< end >>
