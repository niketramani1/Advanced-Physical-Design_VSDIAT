magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1199 -1316 4438 2896
<< locali >>
rect 2583 1443 3160 1477
rect 157 1406 191 1422
rect 1379 1406 1413 1422
rect 191 1372 1379 1406
rect 1413 1372 1662 1406
rect 157 1356 191 1372
rect 1379 1356 1413 1372
rect 77 1298 111 1314
rect 1299 1298 1333 1314
rect 111 1264 1299 1298
rect 1333 1264 1662 1298
rect 77 1248 111 1264
rect 1299 1248 1333 1264
rect 1123 1072 1139 1106
rect 1173 1072 1662 1106
rect 1363 964 1379 998
rect 1413 964 1662 998
rect 2583 893 3160 927
rect 1045 687 1079 703
rect 2583 653 3160 687
rect 1045 637 1079 653
rect 141 603 157 637
rect 191 603 414 637
rect 1203 582 1219 616
rect 1253 582 1662 616
rect 1283 474 1299 508
rect 1333 474 1662 508
rect 1123 282 1139 316
rect 1173 282 1662 316
rect 61 153 77 187
rect 111 153 414 187
rect 1203 174 1219 208
rect 1253 174 1662 208
rect 1045 137 1079 153
rect 2583 103 3160 137
rect 1045 87 1079 103
<< viali >>
rect 157 1372 191 1406
rect 1379 1372 1413 1406
rect 77 1264 111 1298
rect 1299 1264 1333 1298
rect 1139 1072 1173 1106
rect 1379 964 1413 998
rect 1045 653 1079 687
rect 157 603 191 637
rect 1219 582 1253 616
rect 1299 474 1333 508
rect 1139 282 1173 316
rect 77 153 111 187
rect 1219 174 1253 208
rect 1045 103 1079 137
<< metal1 >>
rect 80 1304 108 1500
rect 160 1412 188 1500
rect 145 1406 203 1412
rect 145 1372 157 1406
rect 191 1372 203 1406
rect 145 1366 203 1372
rect 65 1298 123 1304
rect 65 1264 77 1298
rect 111 1264 123 1298
rect 65 1258 123 1264
rect 80 199 108 1258
rect 160 649 188 1366
rect 1142 1118 1170 1500
rect 1133 1106 1179 1118
rect 1133 1072 1139 1106
rect 1173 1072 1179 1106
rect 1133 1060 1179 1072
rect 151 637 197 649
rect 151 603 157 637
rect 191 603 197 637
rect 151 591 197 603
rect 71 187 117 199
rect 71 153 77 187
rect 111 153 117 187
rect 71 141 117 153
rect 80 80 108 141
rect 160 80 188 591
rect 504 421 532 790
rect 900 421 928 790
rect 1030 644 1036 696
rect 1088 644 1094 696
rect 486 369 492 421
rect 544 369 550 421
rect 882 369 888 421
rect 940 369 946 421
rect 504 80 532 369
rect 900 80 928 369
rect 1142 343 1170 1060
rect 1222 738 1250 1500
rect 1302 1310 1330 1500
rect 1382 1418 1410 1500
rect 1373 1412 1419 1418
rect 1367 1406 1425 1412
rect 1367 1372 1379 1406
rect 1413 1372 1425 1406
rect 1367 1366 1425 1372
rect 1373 1360 1419 1366
rect 1293 1304 1339 1310
rect 1287 1298 1345 1304
rect 1287 1264 1299 1298
rect 1333 1264 1345 1298
rect 1287 1258 1345 1264
rect 1293 1252 1339 1258
rect 1210 732 1262 738
rect 1210 674 1262 680
rect 1222 628 1250 674
rect 1213 616 1259 628
rect 1213 582 1219 616
rect 1253 582 1259 616
rect 1213 570 1259 582
rect 1130 337 1182 343
rect 1130 282 1139 285
rect 1173 282 1182 285
rect 1130 279 1182 282
rect 1133 270 1179 279
rect 1030 94 1036 146
rect 1088 94 1094 146
rect 1142 80 1170 270
rect 1222 220 1250 570
rect 1302 520 1330 1252
rect 1382 1010 1410 1360
rect 1788 1218 1836 1610
rect 2212 1218 2262 1612
rect 1780 1166 1786 1218
rect 1838 1166 1844 1218
rect 2205 1166 2211 1218
rect 2263 1166 2269 1218
rect 2602 1211 2630 1580
rect 2998 1211 3026 1580
rect 1373 998 1419 1010
rect 1373 964 1379 998
rect 1413 964 1419 998
rect 1373 952 1419 964
rect 1293 508 1339 520
rect 1293 474 1299 508
rect 1333 474 1339 508
rect 1293 462 1339 474
rect 1213 208 1259 220
rect 1213 174 1219 208
rect 1253 174 1259 208
rect 1213 162 1259 174
rect 1222 80 1250 162
rect 1302 80 1330 462
rect 1382 80 1410 952
rect 1788 428 1836 1166
rect 2212 428 2262 1166
rect 2584 1159 2590 1211
rect 2642 1159 2648 1211
rect 2980 1159 2986 1211
rect 3038 1159 3044 1211
rect 1780 376 1786 428
rect 1838 376 1844 428
rect 2205 376 2211 428
rect 2263 376 2269 428
rect 2602 421 2630 1159
rect 2998 421 3026 1159
rect 1788 80 1836 376
rect 2212 80 2262 376
rect 2584 369 2590 421
rect 2642 369 2648 421
rect 2980 369 2986 421
rect 3038 369 3044 421
rect 2602 80 2630 369
rect 2998 80 3026 369
<< via1 >>
rect 1036 687 1088 696
rect 1036 653 1045 687
rect 1045 653 1079 687
rect 1079 653 1088 687
rect 1036 644 1088 653
rect 492 369 544 421
rect 888 369 940 421
rect 1210 680 1262 732
rect 1130 316 1182 337
rect 1130 285 1139 316
rect 1139 285 1173 316
rect 1173 285 1182 316
rect 1036 137 1088 146
rect 1036 103 1045 137
rect 1045 103 1079 137
rect 1079 103 1088 137
rect 1036 94 1088 103
rect 1786 1166 1838 1218
rect 2211 1166 2263 1218
rect 2590 1159 2642 1211
rect 2986 1159 3038 1211
rect 1786 376 1838 428
rect 2211 376 2263 428
rect 2590 369 2642 421
rect 2986 369 3038 421
<< metal2 >>
rect 1784 1220 1840 1229
rect 1784 1155 1840 1164
rect 2209 1220 2265 1229
rect 2209 1155 2265 1164
rect 2588 1213 2644 1222
rect 2588 1148 2644 1157
rect 2984 1213 3040 1222
rect 2984 1148 3040 1157
rect 1204 720 1210 732
rect 1048 702 1210 720
rect 1036 696 1210 702
rect 1088 692 1210 696
rect 1204 680 1210 692
rect 1262 680 1268 732
rect 1036 638 1088 644
rect 490 423 546 432
rect 490 358 546 367
rect 886 423 942 432
rect 886 358 942 367
rect 1784 430 1840 439
rect 1784 365 1840 374
rect 2209 430 2265 439
rect 2209 365 2265 374
rect 2588 423 2644 432
rect 2588 358 2644 367
rect 2984 423 3040 432
rect 2984 358 3040 367
rect 1124 325 1130 337
rect 1048 297 1130 325
rect 1048 152 1076 297
rect 1124 285 1130 297
rect 1182 285 1188 337
rect 1036 146 1088 152
rect 1036 88 1088 94
<< via2 >>
rect 1784 1218 1840 1220
rect 1784 1166 1786 1218
rect 1786 1166 1838 1218
rect 1838 1166 1840 1218
rect 1784 1164 1840 1166
rect 2209 1218 2265 1220
rect 2209 1166 2211 1218
rect 2211 1166 2263 1218
rect 2263 1166 2265 1218
rect 2209 1164 2265 1166
rect 2588 1211 2644 1213
rect 2588 1159 2590 1211
rect 2590 1159 2642 1211
rect 2642 1159 2644 1211
rect 2588 1157 2644 1159
rect 2984 1211 3040 1213
rect 2984 1159 2986 1211
rect 2986 1159 3038 1211
rect 3038 1159 3040 1211
rect 2984 1157 3040 1159
rect 490 421 546 423
rect 490 369 492 421
rect 492 369 544 421
rect 544 369 546 421
rect 490 367 546 369
rect 886 421 942 423
rect 886 369 888 421
rect 888 369 940 421
rect 940 369 942 421
rect 886 367 942 369
rect 1784 428 1840 430
rect 1784 376 1786 428
rect 1786 376 1838 428
rect 1838 376 1840 428
rect 1784 374 1840 376
rect 2209 428 2265 430
rect 2209 376 2211 428
rect 2211 376 2263 428
rect 2263 376 2265 428
rect 2209 374 2265 376
rect 2588 421 2644 423
rect 2588 369 2590 421
rect 2590 369 2642 421
rect 2642 369 2644 421
rect 2588 367 2644 369
rect 2984 421 3040 423
rect 2984 369 2986 421
rect 2986 369 3038 421
rect 3038 369 3040 421
rect 2984 367 3040 369
<< metal3 >>
rect 1763 1220 1861 1241
rect 1763 1164 1784 1220
rect 1840 1164 1861 1220
rect 1763 1143 1861 1164
rect 2188 1220 2286 1241
rect 2188 1164 2209 1220
rect 2265 1164 2286 1220
rect 2188 1143 2286 1164
rect 2567 1213 2665 1234
rect 2567 1157 2588 1213
rect 2644 1157 2665 1213
rect 2567 1136 2665 1157
rect 2963 1213 3061 1234
rect 2963 1157 2984 1213
rect 3040 1157 3061 1213
rect 2963 1136 3061 1157
rect 469 423 567 444
rect 469 367 490 423
rect 546 367 567 423
rect 469 346 567 367
rect 865 423 963 444
rect 865 367 886 423
rect 942 367 963 423
rect 865 346 963 367
rect 1763 430 1861 451
rect 1763 374 1784 430
rect 1840 374 1861 430
rect 1763 353 1861 374
rect 2188 430 2286 451
rect 2188 374 2209 430
rect 2265 374 2286 430
rect 2188 353 2286 374
rect 2567 423 2665 444
rect 2567 367 2588 423
rect 2644 367 2665 423
rect 2567 346 2665 367
rect 2963 423 3061 444
rect 2963 367 2984 423
rect 3040 367 3061 423
rect 2963 346 3061 367
use pinv_dec  pinv_dec_1
timestamp 1624857261
transform 1 0 320 0 1 0
box 44 0 760 490
use pinv_dec  pinv_dec_0
timestamp 1624857261
transform 1 0 320 0 -1 790
box 44 0 760 490
use contact_17  contact_17_9
timestamp 1624857261
transform 1 0 61 0 1 141
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1624857261
transform 1 0 486 0 1 363
box 0 0 1 1
use contact_7  contact_7_4
timestamp 1624857261
transform 1 0 485 0 1 358
box 0 0 1 1
use contact_17  contact_17_7
timestamp 1624857261
transform 1 0 1123 0 1 270
box 0 0 1 1
use contact_17  contact_17_6
timestamp 1624857261
transform 1 0 1203 0 1 162
box 0 0 1 1
use contact_17  contact_17_5
timestamp 1624857261
transform 1 0 1283 0 1 462
box 0 0 1 1
use contact_14  contact_14_5
timestamp 1624857261
transform 1 0 1033 0 1 87
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1624857261
transform 1 0 1030 0 1 88
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1624857261
transform 1 0 1124 0 1 279
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1624857261
transform 1 0 882 0 1 363
box 0 0 1 1
use contact_7  contact_7_9
timestamp 1624857261
transform 1 0 881 0 1 358
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1624857261
transform 1 0 1779 0 1 365
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1624857261
transform 1 0 1780 0 1 370
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1624857261
transform 1 0 2583 0 1 358
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1624857261
transform 1 0 2584 0 1 363
box 0 0 1 1
use contact_7  contact_7_7
timestamp 1624857261
transform 1 0 2204 0 1 365
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1624857261
transform 1 0 2205 0 1 370
box 0 0 1 1
use contact_7  contact_7_8
timestamp 1624857261
transform 1 0 2979 0 1 358
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1624857261
transform 1 0 2980 0 1 363
box 0 0 1 1
use and2_dec  and2_dec_2
timestamp 1624857261
transform 1 0 1542 0 -1 790
box 70 -56 1636 490
use and2_dec  and2_dec_3
timestamp 1624857261
transform 1 0 1542 0 1 0
box 70 -56 1636 490
use and2_dec  and2_dec_1
timestamp 1624857261
transform 1 0 1542 0 1 790
box 70 -56 1636 490
use contact_17  contact_17_8
timestamp 1624857261
transform 1 0 141 0 1 591
box 0 0 1 1
use contact_17  contact_17_4
timestamp 1624857261
transform 1 0 1203 0 1 570
box 0 0 1 1
use contact_17  contact_17_2
timestamp 1624857261
transform 1 0 1363 0 1 952
box 0 0 1 1
use contact_14  contact_14_4
timestamp 1624857261
transform 1 0 1033 0 1 637
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1624857261
transform 1 0 1030 0 1 638
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1624857261
transform 1 0 1204 0 1 674
box 0 0 1 1
use contact_14  contact_14_3
timestamp 1624857261
transform 1 0 65 0 1 1248
box 0 0 1 1
use contact_17  contact_17_3
timestamp 1624857261
transform 1 0 1123 0 1 1060
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1624857261
transform 1 0 1283 0 1 1252
box 0 0 1 1
use contact_14  contact_14_2
timestamp 1624857261
transform 1 0 1287 0 1 1248
box 0 0 1 1
use contact_19  contact_19_0
timestamp 1624857261
transform 1 0 1780 0 1 1160
box 0 0 1 1
use contact_7  contact_7_0
timestamp 1624857261
transform 1 0 1779 0 1 1155
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1624857261
transform 1 0 2205 0 1 1160
box 0 0 1 1
use contact_7  contact_7_5
timestamp 1624857261
transform 1 0 2204 0 1 1155
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1624857261
transform 1 0 2584 0 1 1153
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1624857261
transform 1 0 2583 0 1 1148
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1624857261
transform 1 0 2980 0 1 1153
box 0 0 1 1
use contact_7  contact_7_6
timestamp 1624857261
transform 1 0 2979 0 1 1148
box 0 0 1 1
use contact_14  contact_14_0
timestamp 1624857261
transform 1 0 1367 0 1 1356
box 0 0 1 1
use contact_14  contact_14_1
timestamp 1624857261
transform 1 0 145 0 1 1356
box 0 0 1 1
use contact_17  contact_17_0
timestamp 1624857261
transform 1 0 1363 0 1 1360
box 0 0 1 1
use and2_dec  and2_dec_0
timestamp 1624857261
transform 1 0 1542 0 -1 1580
box 70 -56 1636 490
<< labels >>
rlabel metal1 s 71 141 117 199 4 in_0
port 1 se
rlabel metal1 s 151 591 197 649 4 in_1
port 2 se
rlabel locali s 2871 120 2871 120 4 out_0
port 3 se
rlabel locali s 2871 670 2871 670 4 out_1
port 4 se
rlabel locali s 2871 910 2871 910 4 out_2
port 5 se
rlabel locali s 2871 1460 2871 1460 4 out_3
port 6 se
rlabel metal3 s 2188 353 2286 451 4 vdd
rlabel metal3 s 865 346 963 444 4 vdd
rlabel metal3 s 2188 1143 2286 1241 4 vdd
rlabel metal3 s 2963 1136 3061 1234 4 vdd
rlabel metal3 s 2963 346 3061 444 4 vdd
port 7 se
rlabel metal3 s 1763 353 1861 451 4 gnd
rlabel metal3 s 469 346 567 444 4 gnd
rlabel metal3 s 2567 346 2665 444 4 gnd
rlabel metal3 s 1763 1143 1861 1241 4 gnd
rlabel metal3 s 2567 1136 2665 1234 4 gnd
port 8 se
<< properties >>
string FIXED_BBOX 0 0 3160 1580
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_END 8767588
string GDS_START 8759764
<< end >>
