magic
tech sky130A
timestamp 1624855461
<< properties >>
string gencell sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield
string parameter m=1
string library sky130
<< end >>
