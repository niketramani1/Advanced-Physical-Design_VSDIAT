magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1288 -1260 1700 2241
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_0
timestamp 1624855509
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_1
timestamp 1624855509
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808520  sky130_fd_pr__dfl1sd__example_55959141808520_0
timestamp 1624855509
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808520  sky130_fd_pr__dfl1sd__example_55959141808520_1
timestamp 1624855509
transform 1 0 412 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 440 981 440 981 0 FreeSans 300 0 0 0 D
flabel comment s 284 981 284 981 0 FreeSans 300 0 0 0 S
flabel comment s 128 981 128 981 0 FreeSans 300 0 0 0 D
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 47461036
string GDS_START 47459082
<< end >>
