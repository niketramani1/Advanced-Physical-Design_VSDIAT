magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1288 -1260 1388 1525
use sky130_fd_pr__hvdfm1sd2__example_55959141808765  sky130_fd_pr__hvdfm1sd2__example_55959141808765_0
timestamp 1624855509
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808765  sky130_fd_pr__hvdfm1sd2__example_55959141808765_1
timestamp 1624855509
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 265 128 265 0 FreeSans 300 0 0 0 D
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 7711776
string GDS_START 7710846
<< end >>
