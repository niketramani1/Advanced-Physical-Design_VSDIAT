magic
tech sky130A
magscale 1 2
timestamp 1624855514
<< nwell >>
rect -83 34302 16087 35388
rect -83 33688 1503 34302
rect 13394 33688 16087 34302
rect -83 33639 16087 33688
rect -83 33296 16088 33639
rect -83 28931 1277 33296
rect 15726 28931 16088 33296
rect -83 28569 16088 28931
rect 9208 27669 16088 27670
rect -83 25726 16088 27669
rect 9388 18442 16134 18626
rect 12530 18340 16134 18442
rect -83 17957 559 18073
rect -83 17290 1195 17957
rect -24 17249 1195 17290
rect -24 17141 1684 17249
rect -24 16925 1699 17141
rect -24 16709 906 16925
rect 15848 16462 16134 18340
rect 9388 16226 16134 16462
rect -143 15554 4963 15840
rect -143 12061 143 15554
rect 15848 14348 16134 16226
rect 12530 14246 16134 14348
rect 9388 14112 16134 14246
rect 15825 12802 16134 14112
rect 14067 12632 16134 12802
rect -143 11797 762 12061
rect -143 11747 2707 11797
rect -143 11629 2092 11747
rect -143 11197 143 11629
rect -143 10911 4703 11197
rect 15825 10003 16134 12632
rect 14067 9717 16134 10003
rect 9783 6446 16090 6804
rect 11655 6075 16090 6446
rect 12966 5550 16090 6075
rect 12966 4209 16090 4662
rect 916 3424 16090 4209
rect -83 726 622 1458
rect 0 -407 12298 293
rect 12806 -29 13078 427
<< pwell >>
rect -32 27756 16032 28480
rect -17 25430 8023 25638
rect 13408 25430 16032 25638
rect -17 24646 16032 25430
rect -17 20277 1121 24646
rect 15599 20277 16032 24646
rect -17 20012 16032 20277
rect -17 18818 1017 20012
rect 7903 19783 16032 20012
rect 10602 19523 16032 19783
rect 15380 19164 16032 19523
rect 7903 18818 16032 19164
rect -17 18814 16032 18818
rect -17 18619 9142 18814
rect -17 18610 9292 18619
rect -17 18206 1834 18610
rect 12875 -357 13215 -207
<< obsli1 >>
rect 0 35322 16000 39534
rect -17 33611 16021 35322
rect -23 28636 16021 33611
rect -23 28624 16000 28636
rect 0 28480 16000 28624
rect -32 27756 16032 28480
rect 0 27623 16000 27756
rect -23 27604 16000 27623
rect -23 25848 16017 27604
rect -17 25792 16017 25848
rect 0 25638 16000 25792
rect -17 25637 16032 25638
rect -23 18814 16032 25637
rect -23 18772 16000 18814
rect -17 18509 16000 18772
rect -17 18206 16017 18509
rect 0 18007 16017 18206
rect -17 17356 16017 18007
rect 0 15714 16017 17356
rect -17 11037 16017 15714
rect 0 9843 16017 11037
rect 0 6738 16000 9843
rect 0 5616 16024 6738
rect 0 4596 16000 5616
rect 0 3490 16024 4596
rect 0 1392 16000 3490
rect -17 792 16000 1392
rect 0 0 16000 792
rect 141 -20 175 0
rect 141 -104 325 -20
rect 418 -97 484 0
rect 141 -300 175 -166
rect 297 -172 331 -166
rect 297 -278 332 -172
rect 518 -269 552 0
rect 694 -239 728 0
rect 766 -16 832 0
rect 870 -269 904 0
rect 1046 -239 1080 0
rect 1222 -269 1256 0
rect 1346 -269 1380 0
rect 1522 -241 1556 0
rect 1698 -269 1732 0
rect 1874 -241 1908 0
rect 2050 -269 2084 0
rect 2123 -11 2189 0
rect 2226 -241 2260 0
rect 2350 -269 2384 0
rect 2526 -241 2560 0
rect 2702 -269 2736 0
rect 2878 -241 2912 0
rect 3054 -269 3088 0
rect 3230 -241 3264 0
rect 3406 -269 3440 0
rect 3582 -241 3616 0
rect 3758 -269 3792 0
rect 3934 -241 3968 0
rect 4110 -269 4144 0
rect 4286 -241 4320 0
rect 4462 -269 4496 0
rect 4638 -241 4672 0
rect 4814 -269 4848 0
rect 4990 -241 5024 0
rect 5166 -269 5200 0
rect 5342 -241 5376 0
rect 5518 -269 5552 0
rect 5694 -241 5728 0
rect 5870 -269 5904 0
rect 5993 -10 6099 0
rect 5994 -241 6028 -10
rect 6170 -269 6204 0
rect 6294 -269 6328 0
rect 6470 -241 6504 0
rect 6646 -269 6680 0
rect 6822 -53 6857 0
rect 6822 -241 6856 -53
rect 7598 -269 7632 0
rect 7774 -241 7808 0
rect 7950 -269 7984 0
rect 8126 -241 8160 0
rect 8250 -269 8284 0
rect 8426 -239 8460 0
rect 8602 -269 8636 0
rect 9058 -82 9092 0
rect 9022 -116 9128 -82
rect 9058 -241 9092 -116
rect 9234 -269 9268 0
rect 9410 -239 9444 0
rect 9586 -269 9620 0
rect 9699 -269 9733 0
rect 9875 -241 9909 0
rect 10051 -269 10085 0
rect 10227 -241 10261 0
rect 10403 -269 10437 0
rect 10528 -241 10562 0
rect 10704 -269 10738 0
rect 10880 -241 10914 0
rect 10950 -43 11016 0
rect 11056 -269 11090 0
rect 11166 -269 11200 0
rect 11342 -241 11376 0
rect 11518 -269 11552 0
rect 11694 -241 11728 0
rect 11804 -269 11838 0
rect 11980 -241 12014 0
rect 12156 -269 12190 0
rect 13658 -19 14001 0
rect 14463 -19 14867 0
rect 13276 -115 13454 -81
rect 13510 -115 13644 -81
rect 13276 -159 13382 -157
rect 13276 -191 13393 -159
rect 297 -300 331 -278
rect 510 -341 12198 -307
rect 12875 -357 13215 -207
rect 13359 -361 13393 -191
rect 13465 -361 13499 -159
rect 13571 -163 13605 -159
rect 13571 -197 13677 -163
rect 13571 -361 13605 -197
<< metal1 >>
rect 12486 -407 12538 -146
<< obsm1 >>
rect 0 35788 16000 39593
rect 0 35373 16004 35788
rect 0 33611 16000 35373
rect -23 25848 16029 33611
rect 0 25637 16000 25848
rect -23 18772 16029 25637
rect 0 18509 16000 18772
rect 0 17889 16012 18509
rect -29 17543 16012 17889
rect 0 15720 16012 17543
rect -23 14179 16012 15720
tri 16012 14179 16023 14190 sw
rect -23 11031 16023 14179
rect 0 9837 16023 11031
rect 0 6738 16000 9837
rect 0 5617 16023 6738
rect 0 4596 16000 5617
rect 0 3490 16023 4596
rect 0 0 16000 3490
rect 52 -26 104 0
tri 203 -26 209 -20 se
rect 209 -26 255 0
tri 181 -48 203 -26 se
rect 203 -40 255 -26
rect 203 -48 247 -40
tri 247 -48 255 -40 nw
tri 135 -94 181 -48 se
rect 135 -293 181 -94
tri 181 -114 247 -48 nw
rect 292 -122 338 0
tri 338 -122 413 -47 sw
rect 428 -51 474 0
rect 776 -16 6111 0
tri 474 -51 508 -17 sw
tri 4551 -22 4557 -16 ne
rect 4557 -22 4685 -16
tri 4685 -22 4691 -16 nw
tri 6766 -51 6817 0 ne
rect 428 -97 3608 -51
tri 3474 -103 3480 -97 ne
rect 3480 -103 3608 -97
rect 4310 -108 5926 -56
rect 5954 -107 6583 -55
rect 6817 -65 6863 0
tri 7114 -17 7131 0 ne
rect 7131 -17 8579 0
tri 8579 -17 8596 0 nw
tri 8661 -17 8678 0 se
rect 8678 -17 9544 0
rect 7092 -97 7624 -45
tri 8608 -70 8661 -17 se
rect 8661 -38 9544 -17
rect 8661 -70 8674 -38
tri 8674 -70 8706 -38 nw
tri 9516 -58 9536 -38 ne
rect 9536 -58 9544 -38
tri 9544 -58 9602 0 sw
tri 10928 -58 10962 -24 se
rect 10962 -58 11008 0
rect 11336 -29 11382 0
tri 9536 -70 9548 -58 ne
rect 9548 -70 11008 -58
rect 7878 -122 8622 -70
tri 8622 -122 8674 -70 nw
rect 9008 -122 9503 -70
tri 9548 -104 9582 -70 ne
rect 9582 -104 11008 -70
rect 292 -150 413 -122
tri 413 -150 441 -122 sw
rect 12486 -146 12538 -24
rect 12736 -119 12976 0
tri 13106 -21 13127 0 ne
rect 292 -353 12239 -150
rect 13127 -169 13155 0
tri 13307 -75 13366 -16 se
rect 13366 -75 13419 0
rect 13264 -121 13419 -75
rect 13471 -75 13499 0
tri 13600 -43 13643 0 ne
tri 13643 -16 13659 0 sw
rect 13643 -43 13659 -16
tri 13499 -75 13531 -43 sw
tri 13643 -59 13659 -43 ne
tri 13659 -59 13702 -16 sw
tri 13659 -74 13674 -59 ne
rect 13471 -121 13631 -75
tri 13155 -169 13183 -141 sw
tri 13246 -169 13264 -151 se
rect 13264 -169 13394 -151
tri 13638 -157 13674 -121 se
rect 13674 -157 13702 -59
rect 13127 -197 13394 -169
rect 13559 -203 13702 -157
rect 12875 -355 13505 -225
tri 15766 -239 15822 -183 se
rect 15822 -239 15874 -167
rect 15051 -295 15874 -239
<< metal2 >>
rect 675 -407 721 488
rect 1084 -407 1130 488
rect 1226 -407 1278 -97
rect 2551 -407 2603 663
rect 3262 -407 3314 57
rect 4471 -407 4523 878
rect 5320 -407 5372 134
rect 5698 -407 5750 407
rect 6150 -407 6202 46
rect 6363 -407 6415 261
rect 7092 -407 7144 -97
rect 7678 -407 7730 211
rect 9049 -407 9101 611
rect 9971 -407 10023 -298
rect 13367 -407 13419 -168
rect 13655 -407 13785 47
rect 15256 -407 15384 4
rect 15522 -407 15574 -170
rect 15741 -407 15781 -164
rect 15943 -407 15983 35167
<< obsm2 >>
rect 42 35223 15983 39593
rect 42 934 15887 35223
rect 42 719 4415 934
rect 42 544 2495 719
rect 42 0 619 544
rect 52 -213 104 0
rect 216 -68 276 0
tri 276 -68 344 0 sw
tri 52 -265 104 -213 ne
tri 104 -223 136 -191 sw
rect 216 -222 344 -68
rect 104 -265 136 -223
tri 104 -295 134 -265 ne
rect 134 -295 136 -265
tri 136 -295 208 -223 sw
tri 134 -347 186 -295 ne
rect 186 -347 432 -295
rect 473 -347 601 0
rect 777 0 1028 544
rect 1186 0 2495 544
tri 1319 -4 1323 0 se
rect 1323 -4 1393 0
tri 1393 -4 1397 0 nw
tri 1245 -78 1319 -4 se
tri 1319 -78 1393 -4 nw
tri 1226 -97 1245 -78 se
rect 1245 -97 1278 -78
tri 1278 -119 1319 -78 nw
rect 1379 -353 2143 -151
rect 2659 113 4415 719
rect 2659 0 3206 113
rect 3370 0 4415 113
tri 3485 -51 3520 -16 se
rect 3520 -51 3572 0
tri 3572 -51 3607 -16 sw
rect 3480 -103 3608 -51
rect 3847 -353 4275 0
tri 4321 -56 4355 -22 se
rect 4355 -56 4407 0
tri 4407 -56 4438 -25 sw
rect 4310 -108 4438 -56
rect 4579 667 15887 934
rect 4579 463 8993 667
rect 4579 190 5642 463
rect 4579 30 5264 190
rect 4557 0 5264 30
rect 4557 -22 4685 0
tri 4701 -108 4809 0 se
rect 4809 -108 5253 0
tri 4659 -150 4701 -108 se
rect 4701 -150 5253 -108
rect 4599 -352 5253 -150
rect 5428 0 5642 190
rect 5806 317 8993 463
rect 5806 102 6307 317
rect 6471 267 8993 317
rect 5806 0 6094 102
tri 5798 -56 5817 -37 se
rect 5817 -56 5870 0
tri 5870 -56 5926 0 sw
rect 5798 -108 5926 -56
rect 5954 -107 6082 0
rect 6258 0 6307 102
rect 6471 144 7622 267
rect 6471 0 7624 144
tri 6455 -33 6471 -17 se
rect 6471 -33 6523 0
rect 6455 -55 6523 -33
tri 6523 -55 6561 -17 sw
rect 6455 -107 6583 -55
rect 6680 -353 6934 0
tri 7065 -27 7092 0 ne
rect 7092 -45 7139 0
tri 7139 -45 7184 0 sw
tri 7496 -45 7541 0 se
rect 7541 -45 7624 0
rect 7092 -97 7220 -45
rect 7496 -97 7624 -45
tri 7144 -137 7184 -97 nw
rect 7786 0 8993 267
tri 7885 -70 7954 -1 se
rect 7954 -70 8006 0
tri 8350 -62 8412 0 se
rect 8412 -62 8424 0
tri 8424 -62 8486 0 nw
rect 7878 -122 8006 -70
tri 8276 -136 8350 -62 se
tri 8350 -136 8424 -62 nw
tri 7730 -180 7769 -141 sw
tri 8232 -180 8276 -136 se
rect 8276 -180 8306 -136
tri 8306 -180 8350 -136 nw
rect 7730 -232 8254 -180
tri 8254 -232 8306 -180 nw
tri 7730 -271 7769 -232 nw
rect 9157 103 15887 667
rect 9157 0 13599 103
rect 13841 60 15887 103
tri 9441 -70 9475 -36 se
rect 9475 -70 9503 0
rect 9879 -33 10033 0
rect 9354 -122 9503 -70
tri 10346 -114 10394 -66 se
rect 10394 -114 10446 0
rect 10505 -8 10831 0
tri 10446 -114 10492 -68 sw
rect 10338 -170 10492 -114
rect 9918 -298 10072 -242
tri 9918 -351 9971 -298 ne
tri 10023 -347 10072 -298 nw
tri 10505 -334 10831 -8 ne
tri 10831 -197 10991 -37 sw
rect 12486 -152 12538 0
rect 12736 -119 12877 0
rect 13308 -168 13472 -112
rect 10831 -334 13040 -197
tri 13308 -227 13367 -168 ne
tri 10831 -347 10844 -334 ne
rect 10844 -347 13040 -334
tri 10844 -351 10848 -347 ne
rect 10848 -351 13040 -347
tri 10848 -353 10850 -351 ne
rect 10850 -353 13040 -351
tri 10850 -357 10854 -353 ne
rect 10854 -357 13040 -353
tri 13419 -221 13472 -168 nw
rect 13841 0 15200 60
rect 15440 4 15887 60
rect 15025 -295 15179 -239
rect 15384 0 15887 4
tri 15384 -82 15466 0 nw
rect 15478 -170 15642 -114
tri 15741 -164 15742 -163 se
rect 15742 -164 15782 0
tri 15482 -210 15522 -170 ne
tri 15574 -232 15636 -170 nw
rect 15781 -181 15782 -164
tri 15781 -182 15782 -181 nw
rect 15822 -295 15874 0
<< metal3 >>
rect 80 -407 204 35290
rect 9173 -407 9239 6954
rect 12564 -407 12778 1534
rect 15716 -407 15782 36548
rect 15848 -407 15914 37505
<< obsm3 >>
rect 80 37585 15914 39593
rect 80 36628 15768 37585
rect 80 35370 15636 36628
rect 284 7034 15636 35370
rect 284 0 9093 7034
rect 283 -218 441 -72
tri 726 -235 736 -225 se
rect 736 -235 802 0
tri 802 -235 882 -155 sw
rect 726 -299 882 -235
rect 1291 -358 2143 0
rect 4527 -357 5527 0
rect 9319 1614 15636 7034
rect 9319 0 12484 1614
rect 9883 -38 10607 0
tri 10607 -38 10645 0 sw
tri 10551 -109 10622 -38 ne
rect 10622 -109 10645 -38
tri 10645 -109 10716 -38 sw
rect 10337 -175 10493 -109
tri 10622 -132 10645 -109 ne
rect 10645 -132 10864 -109
tri 10645 -173 10686 -132 ne
rect 10686 -173 10864 -132
tri 11012 -199 11102 -109 se
rect 11102 -173 11357 -109
tri 11102 -199 11128 -173 nw
tri 10974 -237 11012 -199 se
rect 11012 -237 11041 -199
rect 9922 -260 11041 -237
tri 11041 -260 11102 -199 nw
rect 9922 -301 11000 -260
tri 11000 -301 11041 -260 nw
rect 9922 -303 10068 -301
tri 10068 -303 10070 -301 nw
rect 12858 0 15636 1614
tri 13055 -109 13102 -62 se
rect 13102 -109 13163 0
tri 15332 -83 15415 0 se
rect 15415 -83 15422 0
tri 15422 -83 15505 0 nw
rect 13007 -173 13163 -109
rect 13312 -173 13468 -107
tri 15306 -109 15332 -83 se
rect 15024 -173 15332 -109
tri 15332 -173 15422 -83 nw
rect 15482 -175 15638 -109
rect 15029 -300 15185 -234
<< metal4 >>
rect 0 34750 254 39593
rect 15746 34750 16000 39593
rect 0 13600 254 18593
rect 15746 13600 16000 18593
rect 0 12410 254 13300
rect 15746 12410 16000 13300
rect 0 11240 254 12130
rect 15746 11240 16000 12130
rect 0 10874 522 10940
rect 0 10218 7288 10814
rect 0 9922 254 10158
rect 9418 10874 16000 10940
rect 7752 10218 16000 10814
rect 0 9266 10429 9862
rect 15746 9922 16000 10158
rect 10893 9266 16000 9862
rect 0 9140 522 9206
rect 9418 9140 16000 9206
rect 0 7910 254 8840
rect 15746 7910 16000 8840
rect 0 6940 254 7630
rect 15746 6940 16000 7630
rect 0 5970 254 6660
rect 15746 5970 16000 6660
rect 0 4760 254 5690
rect 15746 4760 16000 5690
rect 0 3550 254 4480
rect 15746 3550 16000 4480
rect 0 2580 193 3270
rect 15794 2580 16000 3270
rect 0 1370 254 2300
rect 15746 1370 16000 2300
rect 0 0 254 1090
rect 15746 0 16000 1090
<< obsm4 >>
rect 334 34670 15666 39593
rect 193 18673 15794 34670
rect 334 13520 15666 18673
rect 193 13380 15794 13520
rect 334 12330 15666 13380
rect 193 12210 15794 12330
rect 334 11160 15666 12210
rect 193 11020 15794 11160
rect 602 10894 9338 11020
rect 7368 10138 7672 10894
rect 334 9942 15666 10138
rect 10509 9286 10813 9942
rect 602 9060 9338 9186
rect 193 8920 15794 9060
rect 334 7830 15666 8920
rect 193 7710 15794 7830
rect 334 6860 15666 7710
rect 193 6740 15794 6860
rect 334 5890 15666 6740
rect 193 5770 15794 5890
rect 334 4680 15666 5770
rect 193 4560 15794 4680
rect 334 3470 15666 4560
rect 193 3350 15794 3470
rect 273 2500 15714 3350
rect 193 2380 15794 2500
rect 334 1290 15666 2380
rect 193 1170 15794 1290
rect 334 0 15666 1170
rect 290 -174 10488 -108
rect 10713 -174 11352 -108
rect 13012 -174 13463 -108
rect 15029 -174 15633 -108
rect 731 -300 15180 -234
<< metal5 >>
rect 2240 20505 14760 32995
rect 0 13600 254 18590
rect 0 12430 254 13280
rect 0 11260 254 12110
rect 0 9140 254 10940
rect 0 7930 254 8820
rect 0 6961 254 7610
rect 0 5990 254 6640
rect 0 4780 254 5670
rect 0 3570 254 4460
rect 15746 13600 16000 18590
rect 15746 12430 16000 13280
rect 15746 11260 16000 12110
rect 15746 9140 16000 10940
rect 15746 7930 16000 8820
rect 15746 6961 16000 7610
rect 15746 5990 16000 6640
rect 15746 4780 16000 5670
rect 15746 3570 16000 4460
rect 0 2600 193 3250
rect 15794 2600 16000 3250
rect 0 1390 254 2280
rect 0 20 254 1070
rect 15746 1390 16000 2280
rect 15746 20 16000 1070
<< obsm5 >>
rect 0 33315 16000 39593
rect 0 20185 1920 33315
rect 15080 20185 16000 33315
rect 0 18910 16000 20185
rect 574 3250 15426 18910
rect 513 2600 15474 3250
rect 574 20 15426 2600
<< labels >>
rlabel metal4 s 0 10218 7288 10814 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel metal4 s 7752 10218 16000 10814 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel metal4 s 0 9266 10429 9862 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel metal4 s 10893 9266 16000 9862 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel metal1 s 12486 -407 12538 -146 8 ANALOG_EN
port 22 nsew signal input
rlabel metal3 s 9173 -407 9239 6954 6 ANALOG_POL
port 26 nsew signal input
rlabel metal2 s 6150 -407 6202 46 8 ANALOG_SEL
port 23 nsew signal input
rlabel metal2 s 5698 -407 5750 407 8 DM[2]
port 6 nsew signal input
rlabel metal2 s 13367 -407 13419 -168 8 DM[1]
port 7 nsew signal input
rlabel metal2 s 9971 -407 10023 -298 8 DM[0]
port 8 nsew signal input
rlabel metal2 s 7092 -407 7144 -97 8 ENABLE_H
port 13 nsew signal input
rlabel metal2 s 7678 -407 7730 211 8 ENABLE_INP_H
port 15 nsew signal input
rlabel metal2 s 2551 -407 2603 663 6 ENABLE_VDDA_H
port 14 nsew signal input
rlabel metal3 s 15716 -407 15782 36548 6 ENABLE_VDDIO
port 24 nsew signal input
rlabel metal2 s 3262 -407 3314 57 8 ENABLE_VSWITCH_H
port 25 nsew signal input
rlabel metal2 s 6363 -407 6415 261 8 HLD_H_N
port 9 nsew signal input
rlabel metal2 s 5320 -407 5372 134 8 HLD_OVR
port 21 nsew signal input
rlabel metal2 s 1084 -407 1130 488 6 IB_MODE_SEL
port 12 nsew signal input
rlabel metal3 s 15848 -407 15914 37505 6 IN
port 10 nsew signal output
rlabel metal3 s 80 -407 204 35290 6 IN_H
port 1 nsew signal output
rlabel metal2 s 9049 -407 9101 611 6 INP_DIS
port 11 nsew signal input
rlabel metal2 s 675 -407 721 488 6 OE_N
port 16 nsew signal input
rlabel metal2 s 4471 -407 4523 878 6 OUT
port 27 nsew signal input
rlabel metal5 s 2240 20505 14760 32995 6 PAD
port 5 nsew signal bidirectional
rlabel metal2 s 15256 -407 15384 4 8 PAD_A_ESD_0_H
port 3 nsew signal bidirectional
rlabel metal2 s 13655 -407 13785 47 8 PAD_A_ESD_1_H
port 4 nsew signal bidirectional
rlabel metal3 s 12564 -407 12778 1534 6 PAD_A_NOESD_H
port 2 nsew signal bidirectional
rlabel metal2 s 15522 -407 15574 -170 8 SLOW
port 19 nsew signal input
rlabel metal2 s 15741 -407 15781 -164 8 TIE_HI_ESD
port 17 nsew signal output
rlabel metal2 s 15943 -407 15983 35167 6 TIE_LO_ESD
port 18 nsew signal output
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 36 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 36 nsew power bidirectional
rlabel metal5 s 15746 1390 16000 2280 6 VCCD
port 36 nsew power bidirectional
rlabel metal4 s 15746 1370 16000 2300 6 VCCD
port 36 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal5 s 15746 20 16000 1070 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal4 s 15746 0 16000 1090 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 31 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 31 nsew power bidirectional
rlabel metal5 s 15794 2600 16000 3250 6 VDDA
port 31 nsew power bidirectional
rlabel metal4 s 15794 2580 16000 3270 6 VDDA
port 31 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 15746 13600 16000 18590 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 15746 3570 16000 4460 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 15746 3550 16000 4480 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 15746 13600 16000 18593 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal5 s 15746 12430 16000 13280 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal4 s 15746 12410 16000 13300 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 9140 522 9206 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 10874 522 10940 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 15746 9140 16000 10940 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 15746 6961 16000 7610 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 15746 9922 16000 10158 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 9418 10874 16000 10940 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 9418 9140 16000 9206 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 15746 6940 16000 7630 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 38 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 38 nsew ground bidirectional
rlabel metal5 s 15746 7930 16000 8820 6 VSSD
port 38 nsew ground bidirectional
rlabel metal4 s 15746 7910 16000 8840 6 VSSD
port 38 nsew ground bidirectional
rlabel metal4 s 0 34750 162 39593 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 15794 34750 16000 39593 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal5 s 15746 4780 16000 5670 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 15746 4760 16000 5690 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 15746 34750 16000 39593 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal5 s 15746 11260 16000 12110 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal4 s 15746 11240 16000 12130 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal5 s 15746 5990 16000 6640 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal4 s 15746 5970 16000 6660 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal2 s 1226 -407 1278 -97 8 VTRIP_SEL
port 20 nsew signal input
<< properties >>
string LEFclass PAD INOUT
string FIXED_BBOX 0 0 16000 39593
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 1807504
string GDS_START 1789672
<< end >>
