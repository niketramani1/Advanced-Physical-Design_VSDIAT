magic
tech sky130A
magscale 1 2
timestamp 1624857261
<< checkpaint >>
rect -1296 -1277 6636 2731
<< nwell >>
rect -36 679 5376 1471
<< locali >>
rect 0 1397 5340 1431
rect 64 636 98 702
rect 915 690 1185 724
rect 196 652 449 686
rect 564 652 817 686
rect 915 669 949 690
rect 1393 674 1769 708
rect 2195 690 2893 724
rect 4073 690 4107 724
rect 0 -17 5340 17
use pinv_19  pinv_19_0
timestamp 1624857261
transform 1 0 2812 0 1 0
box -36 -17 404 1471
use pinv_8  pinv_8_0
timestamp 1624857261
transform 1 0 1688 0 1 0
box -36 -17 836 1471
use pinv_7  pinv_7_0
timestamp 1624857261
transform 1 0 1104 0 1 0
box -36 -17 512 1471
use pinv_0  pinv_0_2
timestamp 1624857261
transform 1 0 0 0 1 0
box -36 -17 404 1471
use pinv_0  pinv_0_1
timestamp 1624857261
transform 1 0 368 0 1 0
box -36 -17 404 1471
use pinv_0  pinv_0_0
timestamp 1624857261
transform 1 0 736 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 4090 707 4090 707 4 Z
port 2 se
rlabel locali s 81 669 81 669 4 A
port 1 se
rlabel locali s 2670 0 2670 0 4 gnd
port 4 se
rlabel locali s 2670 1414 2670 1414 4 vdd
port 3 se
<< properties >>
string FIXED_BBOX 0 0 5340 1414
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_END 8796288
string GDS_START 8794606
<< end >>
