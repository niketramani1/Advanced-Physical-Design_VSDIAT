magic
tech sky130A
magscale 1 2
timestamp 1624855509
<< checkpaint >>
rect -1288 -1260 1584 1323
use sky130_fd_pr__dfl1sd__example_559591418088  sky130_fd_pr__dfl1sd__example_559591418088_0
timestamp 1624855509
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_0
timestamp 1624855509
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808370  sky130_fd_pr__hvdfl1sd__example_55959141808370_0
timestamp 1624855509
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 324 63 324 63 0 FreeSans 300 0 0 0 S
flabel comment s 148 63 148 63 0 FreeSans 300 0 0 0 D
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 639048
string GDS_START 637416
<< end >>
